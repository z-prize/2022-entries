// Copyright Supranational LLC
// Licensed under the Apache License, Version 2.0, see LICENSE-APACHE 
// or the MIT license, see LICENSE-MIT, at your option.
// SPDX-License-Identifier: Apache-2.0 OR MIT

module point_dma
  import config_pkg::*;
  #(
    parameter int ID = 0,
    parameter int C_M00_AXI_ADDR_WIDTH       = 64 ,
    parameter int C_M00_AXI_DATA_WIDTH       = 256,
    parameter int C_M01_AXI_ADDR_WIDTH       = 64 ,
    parameter int C_M01_AXI_DATA_WIDTH       = 256,
    parameter int C_M02_AXI_ADDR_WIDTH       = 64 ,
    parameter int C_M02_AXI_DATA_WIDTH       = 256,
    parameter int C_M03_AXI_ADDR_WIDTH       = 64 ,
    parameter int C_M03_AXI_DATA_WIDTH       = 256,
    parameter int C_M04_AXI_ADDR_WIDTH       = 64 ,
    parameter int C_M04_AXI_DATA_WIDTH       = 256,
    parameter int C_M05_AXI_ADDR_WIDTH       = 64 ,
    parameter int C_M05_AXI_DATA_WIDTH       = 256,
    parameter int C_M06_AXI_ADDR_WIDTH       = 64 ,
    parameter int C_M06_AXI_DATA_WIDTH       = 256,
    parameter int C_M07_AXI_ADDR_WIDTH       = 64 ,
    parameter int C_M07_AXI_DATA_WIDTH       = 256,
    parameter int C_M08_AXI_ADDR_WIDTH       = 64 ,
    parameter int C_M08_AXI_DATA_WIDTH       = 256,
    parameter int C_M09_AXI_ADDR_WIDTH       = 64 ,
    parameter int C_M09_AXI_DATA_WIDTH       = 256,
    parameter int C_M10_AXI_ADDR_WIDTH       = 64 ,
    parameter int C_M10_AXI_DATA_WIDTH       = 256,
    parameter int C_M11_AXI_ADDR_WIDTH       = 64 ,
    parameter int C_M11_AXI_DATA_WIDTH       = 256,
    parameter int C_M12_AXI_ADDR_WIDTH       = 64 ,
    parameter int C_M12_AXI_DATA_WIDTH       = 256,
    parameter int C_M13_AXI_ADDR_WIDTH       = 64 ,
    parameter int C_M13_AXI_DATA_WIDTH       = 256,
    parameter int C_M14_AXI_ADDR_WIDTH       = 64 ,
    parameter int C_M14_AXI_DATA_WIDTH       = 256,
    parameter int C_M15_AXI_ADDR_WIDTH       = 64 ,
    parameter int C_M15_AXI_DATA_WIDTH       = 256,
    parameter int C_M16_AXI_ADDR_WIDTH       = 64 ,
    parameter int C_M16_AXI_DATA_WIDTH       = 256,
    parameter int C_M17_AXI_ADDR_WIDTH       = 64 ,
    parameter int C_M17_AXI_DATA_WIDTH       = 256,
    parameter int C_M18_AXI_ADDR_WIDTH       = 64 ,
    parameter int C_M18_AXI_DATA_WIDTH       = 256,
    parameter int C_M19_AXI_ADDR_WIDTH       = 64 ,
    parameter int C_M19_AXI_DATA_WIDTH       = 256,
    parameter int C_M20_AXI_ADDR_WIDTH       = 64 ,
    parameter int C_M20_AXI_DATA_WIDTH       = 256,
    parameter int C_M21_AXI_ADDR_WIDTH       = 64 ,
    parameter int C_M21_AXI_DATA_WIDTH       = 256,
    parameter int C_M22_AXI_ADDR_WIDTH       = 64 ,
    parameter int C_M22_AXI_DATA_WIDTH       = 256,
    parameter int C_M23_AXI_ADDR_WIDTH       = 64 ,
    parameter int C_M23_AXI_DATA_WIDTH       = 256,
    parameter int C_M24_AXI_ADDR_WIDTH       = 64 ,
    parameter int C_M24_AXI_DATA_WIDTH       = 256,
    parameter int C_M25_AXI_ADDR_WIDTH       = 64 ,
    parameter int C_M25_AXI_DATA_WIDTH       = 256,
    parameter int C_M26_AXI_ADDR_WIDTH       = 64 ,
    parameter int C_M26_AXI_DATA_WIDTH       = 256,
    parameter int C_M27_AXI_ADDR_WIDTH       = 64 ,
    parameter int C_M27_AXI_DATA_WIDTH       = 256,
    parameter int C_M28_AXI_ADDR_WIDTH       = 64 ,
    parameter int C_M28_AXI_DATA_WIDTH       = 256,
    parameter int C_M29_AXI_ADDR_WIDTH       = 64 ,
    parameter int C_M29_AXI_DATA_WIDTH       = 256,
    parameter int C_M30_AXI_ADDR_WIDTH       = 64 ,
    parameter int C_M30_AXI_DATA_WIDTH       = 256,
    parameter int C_M31_AXI_ADDR_WIDTH       = 64 ,
    parameter int C_M31_AXI_DATA_WIDTH       = 256
    )
  (
   input  logic                              clk_i,
   input  logic                              rst_ni,
   input  logic                              start_i,
   output logic                              done_o,

   output logic    [NLANE-1:0][NPPCH-1:0]    re_o,
   input  point_t  [NLANE-1:0][NPPCH-1:0]    rdata_i,
   output fine_t   [NLANE-1:0][NPPCH-1:0]    raddr_o,
   input  coarse_t [NLANE-1:0]               wcoarse_i,
   output coarse_t [NLANE-1:0]               rcoarse_o,

   output logic    [NLANE-1:0][NPPCH-1:0]    we_o,
   output point_t  [NLANE-1:0][NPPCH-1:0]    wdata_o,
   output fine_t   [NLANE-1:0][NPPCH-1:0]    waddr_o,
   output coarse_t [NLANE-1:0]               wcoarse_o,
   input  coarse_t [NLANE-1:0]               rcoarse_i,

   output 				     beat_id_t dbg_ch0_wbeat,
   output 				     beat_id_t dbg_ch0_rbeat,
   output 				     beat_id_t dbg_ch8_wbeat,
   output 				     beat_id_t dbg_ch8_rbeat,
   output logic [15:0]			     dbg_wstep,
   output logic [15:0]			     dbg_rstep,

   // Tool generated ports.
   output logic                              m00_axi_awvalid,
   input  logic                              m00_axi_awready,
   output logic [C_M00_AXI_ADDR_WIDTH-1:0]   m00_axi_awaddr ,
   output logic [8-1:0]                      m00_axi_awlen  ,
   output logic                              m00_axi_wvalid ,
   input  logic                              m00_axi_wready ,
   output logic [C_M00_AXI_DATA_WIDTH-1:0]   m00_axi_wdata  ,
   output logic [C_M00_AXI_DATA_WIDTH/8-1:0] m00_axi_wstrb  ,
   output logic                              m00_axi_wlast  ,
   input  logic                              m00_axi_bvalid ,
   output logic                              m00_axi_bready ,
   output logic                              m00_axi_arvalid,
   input  logic                              m00_axi_arready,
   output logic [C_M00_AXI_ADDR_WIDTH-1:0]   m00_axi_araddr ,
   output logic [8-1:0]                      m00_axi_arlen  ,
   input  logic                              m00_axi_rvalid ,
   output logic                              m00_axi_rready ,
   input  logic [C_M00_AXI_DATA_WIDTH-1:0]   m00_axi_rdata  ,
   input  logic                              m00_axi_rlast  ,

   output logic                              m01_axi_awvalid,
   input  logic                              m01_axi_awready,
   output logic [C_M01_AXI_ADDR_WIDTH-1:0]   m01_axi_awaddr ,
   output logic [8-1:0]                      m01_axi_awlen  ,
   output logic                              m01_axi_wvalid ,
   input  logic                              m01_axi_wready ,
   output logic [C_M01_AXI_DATA_WIDTH-1:0]   m01_axi_wdata  ,
   output logic [C_M01_AXI_DATA_WIDTH/8-1:0] m01_axi_wstrb  ,
   output logic                              m01_axi_wlast  ,
   input  logic                              m01_axi_bvalid ,
   output logic                              m01_axi_bready ,
   output logic                              m01_axi_arvalid,
   input  logic                              m01_axi_arready,
   output logic [C_M01_AXI_ADDR_WIDTH-1:0]   m01_axi_araddr ,
   output logic [8-1:0]                      m01_axi_arlen  ,
   input  logic                              m01_axi_rvalid ,
   output logic                              m01_axi_rready ,
   input  logic [C_M01_AXI_DATA_WIDTH-1:0]   m01_axi_rdata  ,
   input  logic                              m01_axi_rlast  ,

   output logic                              m02_axi_awvalid,
   input  logic                              m02_axi_awready,
   output logic [C_M02_AXI_ADDR_WIDTH-1:0]   m02_axi_awaddr ,
   output logic [8-1:0]                      m02_axi_awlen  ,
   output logic                              m02_axi_wvalid ,
   input  logic                              m02_axi_wready ,
   output logic [C_M02_AXI_DATA_WIDTH-1:0]   m02_axi_wdata  ,
   output logic [C_M02_AXI_DATA_WIDTH/8-1:0] m02_axi_wstrb  ,
   output logic                              m02_axi_wlast  ,
   input  logic                              m02_axi_bvalid ,
   output logic                              m02_axi_bready ,
   output logic                              m02_axi_arvalid,
   input  logic                              m02_axi_arready,
   output logic [C_M02_AXI_ADDR_WIDTH-1:0]   m02_axi_araddr ,
   output logic [8-1:0]                      m02_axi_arlen  ,
   input  logic                              m02_axi_rvalid ,
   output logic                              m02_axi_rready ,
   input  logic [C_M02_AXI_DATA_WIDTH-1:0]   m02_axi_rdata  ,
   input  logic                              m02_axi_rlast  ,

   output logic                              m03_axi_awvalid,
   input  logic                              m03_axi_awready,
   output logic [C_M03_AXI_ADDR_WIDTH-1:0]   m03_axi_awaddr ,
   output logic [8-1:0]                      m03_axi_awlen  ,
   output logic                              m03_axi_wvalid ,
   input  logic                              m03_axi_wready ,
   output logic [C_M03_AXI_DATA_WIDTH-1:0]   m03_axi_wdata  ,
   output logic [C_M03_AXI_DATA_WIDTH/8-1:0] m03_axi_wstrb  ,
   output logic                              m03_axi_wlast  ,
   input  logic                              m03_axi_bvalid ,
   output logic                              m03_axi_bready ,
   output logic                              m03_axi_arvalid,
   input  logic                              m03_axi_arready,
   output logic [C_M03_AXI_ADDR_WIDTH-1:0]   m03_axi_araddr ,
   output logic [8-1:0]                      m03_axi_arlen  ,
   input  logic                              m03_axi_rvalid ,
   output logic                              m03_axi_rready ,
   input  logic [C_M03_AXI_DATA_WIDTH-1:0]   m03_axi_rdata  ,
   input  logic                              m03_axi_rlast  ,

   output logic                              m04_axi_awvalid,
   input  logic                              m04_axi_awready,
   output logic [C_M04_AXI_ADDR_WIDTH-1:0]   m04_axi_awaddr ,
   output logic [8-1:0]                      m04_axi_awlen  ,
   output logic                              m04_axi_wvalid ,
   input  logic                              m04_axi_wready ,
   output logic [C_M04_AXI_DATA_WIDTH-1:0]   m04_axi_wdata  ,
   output logic [C_M04_AXI_DATA_WIDTH/8-1:0] m04_axi_wstrb  ,
   output logic                              m04_axi_wlast  ,
   input  logic                              m04_axi_bvalid ,
   output logic                              m04_axi_bready ,
   output logic                              m04_axi_arvalid,
   input  logic                              m04_axi_arready,
   output logic [C_M04_AXI_ADDR_WIDTH-1:0]   m04_axi_araddr ,
   output logic [8-1:0]                      m04_axi_arlen  ,
   input  logic                              m04_axi_rvalid ,
   output logic                              m04_axi_rready ,
   input  logic [C_M04_AXI_DATA_WIDTH-1:0]   m04_axi_rdata  ,
   input  logic                              m04_axi_rlast  ,

   output logic                              m05_axi_awvalid,
   input  logic                              m05_axi_awready,
   output logic [C_M05_AXI_ADDR_WIDTH-1:0]   m05_axi_awaddr ,
   output logic [8-1:0]                      m05_axi_awlen  ,
   output logic                              m05_axi_wvalid ,
   input  logic                              m05_axi_wready ,
   output logic [C_M05_AXI_DATA_WIDTH-1:0]   m05_axi_wdata  ,
   output logic [C_M05_AXI_DATA_WIDTH/8-1:0] m05_axi_wstrb  ,
   output logic                              m05_axi_wlast  ,
   input  logic                              m05_axi_bvalid ,
   output logic                              m05_axi_bready ,
   output logic                              m05_axi_arvalid,
   input  logic                              m05_axi_arready,
   output logic [C_M05_AXI_ADDR_WIDTH-1:0]   m05_axi_araddr ,
   output logic [8-1:0]                      m05_axi_arlen  ,
   input  logic                              m05_axi_rvalid ,
   output logic                              m05_axi_rready ,
   input  logic [C_M05_AXI_DATA_WIDTH-1:0]   m05_axi_rdata  ,
   input  logic                              m05_axi_rlast  ,

   output logic                              m06_axi_awvalid,
   input  logic                              m06_axi_awready,
   output logic [C_M06_AXI_ADDR_WIDTH-1:0]   m06_axi_awaddr ,
   output logic [8-1:0]                      m06_axi_awlen  ,
   output logic                              m06_axi_wvalid ,
   input  logic                              m06_axi_wready ,
   output logic [C_M06_AXI_DATA_WIDTH-1:0]   m06_axi_wdata  ,
   output logic [C_M06_AXI_DATA_WIDTH/8-1:0] m06_axi_wstrb  ,
   output logic                              m06_axi_wlast  ,
   input  logic                              m06_axi_bvalid ,
   output logic                              m06_axi_bready ,
   output logic                              m06_axi_arvalid,
   input  logic                              m06_axi_arready,
   output logic [C_M06_AXI_ADDR_WIDTH-1:0]   m06_axi_araddr ,
   output logic [8-1:0]                      m06_axi_arlen  ,
   input  logic                              m06_axi_rvalid ,
   output logic                              m06_axi_rready ,
   input  logic [C_M06_AXI_DATA_WIDTH-1:0]   m06_axi_rdata  ,
   input  logic                              m06_axi_rlast  ,

   output logic                              m07_axi_awvalid,
   input  logic                              m07_axi_awready,
   output logic [C_M07_AXI_ADDR_WIDTH-1:0]   m07_axi_awaddr ,
   output logic [8-1:0]                      m07_axi_awlen  ,
   output logic                              m07_axi_wvalid ,
   input  logic                              m07_axi_wready ,
   output logic [C_M07_AXI_DATA_WIDTH-1:0]   m07_axi_wdata  ,
   output logic [C_M07_AXI_DATA_WIDTH/8-1:0] m07_axi_wstrb  ,
   output logic                              m07_axi_wlast  ,
   input  logic                              m07_axi_bvalid ,
   output logic                              m07_axi_bready ,
   output logic                              m07_axi_arvalid,
   input  logic                              m07_axi_arready,
   output logic [C_M07_AXI_ADDR_WIDTH-1:0]   m07_axi_araddr ,
   output logic [8-1:0]                      m07_axi_arlen  ,
   input  logic                              m07_axi_rvalid ,
   output logic                              m07_axi_rready ,
   input  logic [C_M07_AXI_DATA_WIDTH-1:0]   m07_axi_rdata  ,
   input  logic                              m07_axi_rlast  ,

   output logic                              m08_axi_awvalid,
   input  logic                              m08_axi_awready,
   output logic [C_M08_AXI_ADDR_WIDTH-1:0]   m08_axi_awaddr ,
   output logic [8-1:0]                      m08_axi_awlen  ,
   output logic                              m08_axi_wvalid ,
   input  logic                              m08_axi_wready ,
   output logic [C_M08_AXI_DATA_WIDTH-1:0]   m08_axi_wdata  ,
   output logic [C_M08_AXI_DATA_WIDTH/8-1:0] m08_axi_wstrb  ,
   output logic                              m08_axi_wlast  ,
   input  logic                              m08_axi_bvalid ,
   output logic                              m08_axi_bready ,
   output logic                              m08_axi_arvalid,
   input  logic                              m08_axi_arready,
   output logic [C_M08_AXI_ADDR_WIDTH-1:0]   m08_axi_araddr ,
   output logic [8-1:0]                      m08_axi_arlen  ,
   input  logic                              m08_axi_rvalid ,
   output logic                              m08_axi_rready ,
   input  logic [C_M08_AXI_DATA_WIDTH-1:0]   m08_axi_rdata  ,
   input  logic                              m08_axi_rlast  ,

   output logic                              m09_axi_awvalid,
   input  logic                              m09_axi_awready,
   output logic [C_M09_AXI_ADDR_WIDTH-1:0]   m09_axi_awaddr ,
   output logic [8-1:0]                      m09_axi_awlen  ,
   output logic                              m09_axi_wvalid ,
   input  logic                              m09_axi_wready ,
   output logic [C_M09_AXI_DATA_WIDTH-1:0]   m09_axi_wdata  ,
   output logic [C_M09_AXI_DATA_WIDTH/8-1:0] m09_axi_wstrb  ,
   output logic                              m09_axi_wlast  ,
   input  logic                              m09_axi_bvalid ,
   output logic                              m09_axi_bready ,
   output logic                              m09_axi_arvalid,
   input  logic                              m09_axi_arready,
   output logic [C_M09_AXI_ADDR_WIDTH-1:0]   m09_axi_araddr ,
   output logic [8-1:0]                      m09_axi_arlen  ,
   input  logic                              m09_axi_rvalid ,
   output logic                              m09_axi_rready ,
   input  logic [C_M09_AXI_DATA_WIDTH-1:0]   m09_axi_rdata  ,
   input  logic                              m09_axi_rlast  ,

   output logic                              m10_axi_awvalid,
   input  logic                              m10_axi_awready,
   output logic [C_M10_AXI_ADDR_WIDTH-1:0]   m10_axi_awaddr ,
   output logic [8-1:0]                      m10_axi_awlen  ,
   output logic                              m10_axi_wvalid ,
   input  logic                              m10_axi_wready ,
   output logic [C_M10_AXI_DATA_WIDTH-1:0]   m10_axi_wdata  ,
   output logic [C_M10_AXI_DATA_WIDTH/8-1:0] m10_axi_wstrb  ,
   output logic                              m10_axi_wlast  ,
   input  logic                              m10_axi_bvalid ,
   output logic                              m10_axi_bready ,
   output logic                              m10_axi_arvalid,
   input  logic                              m10_axi_arready,
   output logic [C_M10_AXI_ADDR_WIDTH-1:0]   m10_axi_araddr ,
   output logic [8-1:0]                      m10_axi_arlen  ,
   input  logic                              m10_axi_rvalid ,
   output logic                              m10_axi_rready ,
   input  logic [C_M10_AXI_DATA_WIDTH-1:0]   m10_axi_rdata  ,
   input  logic                              m10_axi_rlast  ,

   output logic                              m11_axi_awvalid,
   input  logic                              m11_axi_awready,
   output logic [C_M11_AXI_ADDR_WIDTH-1:0]   m11_axi_awaddr ,
   output logic [8-1:0]                      m11_axi_awlen  ,
   output logic                              m11_axi_wvalid ,
   input  logic                              m11_axi_wready ,
   output logic [C_M11_AXI_DATA_WIDTH-1:0]   m11_axi_wdata  ,
   output logic [C_M11_AXI_DATA_WIDTH/8-1:0] m11_axi_wstrb  ,
   output logic                              m11_axi_wlast  ,
   input  logic                              m11_axi_bvalid ,
   output logic                              m11_axi_bready ,
   output logic                              m11_axi_arvalid,
   input  logic                              m11_axi_arready,
   output logic [C_M11_AXI_ADDR_WIDTH-1:0]   m11_axi_araddr ,
   output logic [8-1:0]                      m11_axi_arlen  ,
   input  logic                              m11_axi_rvalid ,
   output logic                              m11_axi_rready ,
   input  logic [C_M11_AXI_DATA_WIDTH-1:0]   m11_axi_rdata  ,
   input  logic                              m11_axi_rlast  ,

   output logic                              m12_axi_awvalid,
   input  logic                              m12_axi_awready,
   output logic [C_M12_AXI_ADDR_WIDTH-1:0]   m12_axi_awaddr ,
   output logic [8-1:0]                      m12_axi_awlen  ,
   output logic                              m12_axi_wvalid ,
   input  logic                              m12_axi_wready ,
   output logic [C_M12_AXI_DATA_WIDTH-1:0]   m12_axi_wdata  ,
   output logic [C_M12_AXI_DATA_WIDTH/8-1:0] m12_axi_wstrb  ,
   output logic                              m12_axi_wlast  ,
   input  logic                              m12_axi_bvalid ,
   output logic                              m12_axi_bready ,
   output logic                              m12_axi_arvalid,
   input  logic                              m12_axi_arready,
   output logic [C_M12_AXI_ADDR_WIDTH-1:0]   m12_axi_araddr ,
   output logic [8-1:0]                      m12_axi_arlen  ,
   input  logic                              m12_axi_rvalid ,
   output logic                              m12_axi_rready ,
   input  logic [C_M12_AXI_DATA_WIDTH-1:0]   m12_axi_rdata  ,
   input  logic                              m12_axi_rlast  ,

   output logic                              m13_axi_awvalid,
   input  logic                              m13_axi_awready,
   output logic [C_M13_AXI_ADDR_WIDTH-1:0]   m13_axi_awaddr ,
   output logic [8-1:0]                      m13_axi_awlen  ,
   output logic                              m13_axi_wvalid ,
   input  logic                              m13_axi_wready ,
   output logic [C_M13_AXI_DATA_WIDTH-1:0]   m13_axi_wdata  ,
   output logic [C_M13_AXI_DATA_WIDTH/8-1:0] m13_axi_wstrb  ,
   output logic                              m13_axi_wlast  ,
   input  logic                              m13_axi_bvalid ,
   output logic                              m13_axi_bready ,
   output logic                              m13_axi_arvalid,
   input  logic                              m13_axi_arready,
   output logic [C_M13_AXI_ADDR_WIDTH-1:0]   m13_axi_araddr ,
   output logic [8-1:0]                      m13_axi_arlen  ,
   input  logic                              m13_axi_rvalid ,
   output logic                              m13_axi_rready ,
   input  logic [C_M13_AXI_DATA_WIDTH-1:0]   m13_axi_rdata  ,
   input  logic                              m13_axi_rlast  ,

   output logic                              m14_axi_awvalid,
   input  logic                              m14_axi_awready,
   output logic [C_M14_AXI_ADDR_WIDTH-1:0]   m14_axi_awaddr ,
   output logic [8-1:0]                      m14_axi_awlen  ,
   output logic                              m14_axi_wvalid ,
   input  logic                              m14_axi_wready ,
   output logic [C_M14_AXI_DATA_WIDTH-1:0]   m14_axi_wdata  ,
   output logic [C_M14_AXI_DATA_WIDTH/8-1:0] m14_axi_wstrb  ,
   output logic                              m14_axi_wlast  ,
   input  logic                              m14_axi_bvalid ,
   output logic                              m14_axi_bready ,
   output logic                              m14_axi_arvalid,
   input  logic                              m14_axi_arready,
   output logic [C_M14_AXI_ADDR_WIDTH-1:0]   m14_axi_araddr ,
   output logic [8-1:0]                      m14_axi_arlen  ,
   input  logic                              m14_axi_rvalid ,
   output logic                              m14_axi_rready ,
   input  logic [C_M14_AXI_DATA_WIDTH-1:0]   m14_axi_rdata  ,
   input  logic                              m14_axi_rlast  ,

   output logic                              m15_axi_awvalid,
   input  logic                              m15_axi_awready,
   output logic [C_M15_AXI_ADDR_WIDTH-1:0]   m15_axi_awaddr ,
   output logic [8-1:0]                      m15_axi_awlen  ,
   output logic                              m15_axi_wvalid ,
   input  logic                              m15_axi_wready ,
   output logic [C_M15_AXI_DATA_WIDTH-1:0]   m15_axi_wdata  ,
   output logic [C_M15_AXI_DATA_WIDTH/8-1:0] m15_axi_wstrb  ,
   output logic                              m15_axi_wlast  ,
   input  logic                              m15_axi_bvalid ,
   output logic                              m15_axi_bready ,
   output logic                              m15_axi_arvalid,
   input  logic                              m15_axi_arready,
   output logic [C_M15_AXI_ADDR_WIDTH-1:0]   m15_axi_araddr ,
   output logic [8-1:0]                      m15_axi_arlen  ,
   input  logic                              m15_axi_rvalid ,
   output logic                              m15_axi_rready ,
   input  logic [C_M15_AXI_DATA_WIDTH-1:0]   m15_axi_rdata  ,
   input  logic                              m15_axi_rlast  ,

   output logic                              m16_axi_awvalid,
   input  logic                              m16_axi_awready,
   output logic [C_M06_AXI_ADDR_WIDTH-1:0]   m16_axi_awaddr ,
   output logic [8-1:0]                      m16_axi_awlen  ,
   output logic                              m16_axi_wvalid ,
   input  logic                              m16_axi_wready ,
   output logic [C_M06_AXI_DATA_WIDTH-1:0]   m16_axi_wdata  ,
   output logic [C_M06_AXI_DATA_WIDTH/8-1:0] m16_axi_wstrb  ,
   output logic                              m16_axi_wlast  ,
   input  logic                              m16_axi_bvalid ,
   output logic                              m16_axi_bready ,
   output logic                              m16_axi_arvalid,
   input  logic                              m16_axi_arready,
   output logic [C_M06_AXI_ADDR_WIDTH-1:0]   m16_axi_araddr ,
   output logic [8-1:0]                      m16_axi_arlen  ,
   input  logic                              m16_axi_rvalid ,
   output logic                              m16_axi_rready ,
   input  logic [C_M06_AXI_DATA_WIDTH-1:0]   m16_axi_rdata  ,
   input  logic                              m16_axi_rlast  ,

   output logic                              m17_axi_awvalid,
   input  logic                              m17_axi_awready,
   output logic [C_M07_AXI_ADDR_WIDTH-1:0]   m17_axi_awaddr ,
   output logic [8-1:0]                      m17_axi_awlen  ,
   output logic                              m17_axi_wvalid ,
   input  logic                              m17_axi_wready ,
   output logic [C_M07_AXI_DATA_WIDTH-1:0]   m17_axi_wdata  ,
   output logic [C_M07_AXI_DATA_WIDTH/8-1:0] m17_axi_wstrb  ,
   output logic                              m17_axi_wlast  ,
   input  logic                              m17_axi_bvalid ,
   output logic                              m17_axi_bready ,
   output logic                              m17_axi_arvalid,
   input  logic                              m17_axi_arready,
   output logic [C_M07_AXI_ADDR_WIDTH-1:0]   m17_axi_araddr ,
   output logic [8-1:0]                      m17_axi_arlen  ,
   input  logic                              m17_axi_rvalid ,
   output logic                              m17_axi_rready ,
   input  logic [C_M07_AXI_DATA_WIDTH-1:0]   m17_axi_rdata  ,
   input  logic                              m17_axi_rlast  ,

   output logic                              m18_axi_awvalid,
   input  logic                              m18_axi_awready,
   output logic [C_M08_AXI_ADDR_WIDTH-1:0]   m18_axi_awaddr ,
   output logic [8-1:0]                      m18_axi_awlen  ,
   output logic                              m18_axi_wvalid ,
   input  logic                              m18_axi_wready ,
   output logic [C_M08_AXI_DATA_WIDTH-1:0]   m18_axi_wdata  ,
   output logic [C_M08_AXI_DATA_WIDTH/8-1:0] m18_axi_wstrb  ,
   output logic                              m18_axi_wlast  ,
   input  logic                              m18_axi_bvalid ,
   output logic                              m18_axi_bready ,
   output logic                              m18_axi_arvalid,
   input  logic                              m18_axi_arready,
   output logic [C_M08_AXI_ADDR_WIDTH-1:0]   m18_axi_araddr ,
   output logic [8-1:0]                      m18_axi_arlen  ,
   input  logic                              m18_axi_rvalid ,
   output logic                              m18_axi_rready ,
   input  logic [C_M08_AXI_DATA_WIDTH-1:0]   m18_axi_rdata  ,
   input  logic                              m18_axi_rlast  ,

   output logic                              m19_axi_awvalid,
   input  logic                              m19_axi_awready,
   output logic [C_M09_AXI_ADDR_WIDTH-1:0]   m19_axi_awaddr ,
   output logic [8-1:0]                      m19_axi_awlen  ,
   output logic                              m19_axi_wvalid ,
   input  logic                              m19_axi_wready ,
   output logic [C_M09_AXI_DATA_WIDTH-1:0]   m19_axi_wdata  ,
   output logic [C_M09_AXI_DATA_WIDTH/8-1:0] m19_axi_wstrb  ,
   output logic                              m19_axi_wlast  ,
   input  logic                              m19_axi_bvalid ,
   output logic                              m19_axi_bready ,
   output logic                              m19_axi_arvalid,
   input  logic                              m19_axi_arready,
   output logic [C_M09_AXI_ADDR_WIDTH-1:0]   m19_axi_araddr ,
   output logic [8-1:0]                      m19_axi_arlen  ,
   input  logic                              m19_axi_rvalid ,
   output logic                              m19_axi_rready ,
   input  logic [C_M09_AXI_DATA_WIDTH-1:0]   m19_axi_rdata  ,
   input  logic                              m19_axi_rlast  ,

   output logic                              m20_axi_awvalid,
   input  logic                              m20_axi_awready,
   output logic [C_M10_AXI_ADDR_WIDTH-1:0]   m20_axi_awaddr ,
   output logic [8-1:0]                      m20_axi_awlen  ,
   output logic                              m20_axi_wvalid ,
   input  logic                              m20_axi_wready ,
   output logic [C_M10_AXI_DATA_WIDTH-1:0]   m20_axi_wdata  ,
   output logic [C_M10_AXI_DATA_WIDTH/8-1:0] m20_axi_wstrb  ,
   output logic                              m20_axi_wlast  ,
   input  logic                              m20_axi_bvalid ,
   output logic                              m20_axi_bready ,
   output logic                              m20_axi_arvalid,
   input  logic                              m20_axi_arready,
   output logic [C_M10_AXI_ADDR_WIDTH-1:0]   m20_axi_araddr ,
   output logic [8-1:0]                      m20_axi_arlen  ,
   input  logic                              m20_axi_rvalid ,
   output logic                              m20_axi_rready ,
   input  logic [C_M10_AXI_DATA_WIDTH-1:0]   m20_axi_rdata  ,
   input  logic                              m20_axi_rlast  ,

   output logic                              m21_axi_awvalid,
   input  logic                              m21_axi_awready,
   output logic [C_M11_AXI_ADDR_WIDTH-1:0]   m21_axi_awaddr ,
   output logic [8-1:0]                      m21_axi_awlen  ,
   output logic                              m21_axi_wvalid ,
   input  logic                              m21_axi_wready ,
   output logic [C_M11_AXI_DATA_WIDTH-1:0]   m21_axi_wdata  ,
   output logic [C_M11_AXI_DATA_WIDTH/8-1:0] m21_axi_wstrb  ,
   output logic                              m21_axi_wlast  ,
   input  logic                              m21_axi_bvalid ,
   output logic                              m21_axi_bready ,
   output logic                              m21_axi_arvalid,
   input  logic                              m21_axi_arready,
   output logic [C_M11_AXI_ADDR_WIDTH-1:0]   m21_axi_araddr ,
   output logic [8-1:0]                      m21_axi_arlen  ,
   input  logic                              m21_axi_rvalid ,
   output logic                              m21_axi_rready ,
   input  logic [C_M11_AXI_DATA_WIDTH-1:0]   m21_axi_rdata  ,
   input  logic                              m21_axi_rlast  ,

   output logic                              m22_axi_awvalid,
   input  logic                              m22_axi_awready,
   output logic [C_M02_AXI_ADDR_WIDTH-1:0]   m22_axi_awaddr ,
   output logic [8-1:0]                      m22_axi_awlen  ,
   output logic                              m22_axi_wvalid ,
   input  logic                              m22_axi_wready ,
   output logic [C_M02_AXI_DATA_WIDTH-1:0]   m22_axi_wdata  ,
   output logic [C_M02_AXI_DATA_WIDTH/8-1:0] m22_axi_wstrb  ,
   output logic                              m22_axi_wlast  ,
   input  logic                              m22_axi_bvalid ,
   output logic                              m22_axi_bready ,
   output logic                              m22_axi_arvalid,
   input  logic                              m22_axi_arready,
   output logic [C_M02_AXI_ADDR_WIDTH-1:0]   m22_axi_araddr ,
   output logic [8-1:0]                      m22_axi_arlen  ,
   input  logic                              m22_axi_rvalid ,
   output logic                              m22_axi_rready ,
   input  logic [C_M02_AXI_DATA_WIDTH-1:0]   m22_axi_rdata  ,
   input  logic                              m22_axi_rlast  ,

   output logic                              m23_axi_awvalid,
   input  logic                              m23_axi_awready,
   output logic [C_M03_AXI_ADDR_WIDTH-1:0]   m23_axi_awaddr ,
   output logic [8-1:0]                      m23_axi_awlen  ,
   output logic                              m23_axi_wvalid ,
   input  logic                              m23_axi_wready ,
   output logic [C_M03_AXI_DATA_WIDTH-1:0]   m23_axi_wdata  ,
   output logic [C_M03_AXI_DATA_WIDTH/8-1:0] m23_axi_wstrb  ,
   output logic                              m23_axi_wlast  ,
   input  logic                              m23_axi_bvalid ,
   output logic                              m23_axi_bready ,
   output logic                              m23_axi_arvalid,
   input  logic                              m23_axi_arready,
   output logic [C_M03_AXI_ADDR_WIDTH-1:0]   m23_axi_araddr ,
   output logic [8-1:0]                      m23_axi_arlen  ,
   input  logic                              m23_axi_rvalid ,
   output logic                              m23_axi_rready ,
   input  logic [C_M03_AXI_DATA_WIDTH-1:0]   m23_axi_rdata  ,
   input  logic                              m23_axi_rlast  ,

   output logic                              m24_axi_awvalid,
   input  logic                              m24_axi_awready,
   output logic [C_M04_AXI_ADDR_WIDTH-1:0]   m24_axi_awaddr ,
   output logic [8-1:0]                      m24_axi_awlen  ,
   output logic                              m24_axi_wvalid ,
   input  logic                              m24_axi_wready ,
   output logic [C_M04_AXI_DATA_WIDTH-1:0]   m24_axi_wdata  ,
   output logic [C_M04_AXI_DATA_WIDTH/8-1:0] m24_axi_wstrb  ,
   output logic                              m24_axi_wlast  ,
   input  logic                              m24_axi_bvalid ,
   output logic                              m24_axi_bready ,
   output logic                              m24_axi_arvalid,
   input  logic                              m24_axi_arready,
   output logic [C_M04_AXI_ADDR_WIDTH-1:0]   m24_axi_araddr ,
   output logic [8-1:0]                      m24_axi_arlen  ,
   input  logic                              m24_axi_rvalid ,
   output logic                              m24_axi_rready ,
   input  logic [C_M04_AXI_DATA_WIDTH-1:0]   m24_axi_rdata  ,
   input  logic                              m24_axi_rlast  ,

   output logic                              m25_axi_awvalid,
   input  logic                              m25_axi_awready,
   output logic [C_M05_AXI_ADDR_WIDTH-1:0]   m25_axi_awaddr ,
   output logic [8-1:0]                      m25_axi_awlen  ,
   output logic                              m25_axi_wvalid ,
   input  logic                              m25_axi_wready ,
   output logic [C_M05_AXI_DATA_WIDTH-1:0]   m25_axi_wdata  ,
   output logic [C_M05_AXI_DATA_WIDTH/8-1:0] m25_axi_wstrb  ,
   output logic                              m25_axi_wlast  ,
   input  logic                              m25_axi_bvalid ,
   output logic                              m25_axi_bready ,
   output logic                              m25_axi_arvalid,
   input  logic                              m25_axi_arready,
   output logic [C_M05_AXI_ADDR_WIDTH-1:0]   m25_axi_araddr ,
   output logic [8-1:0]                      m25_axi_arlen  ,
   input  logic                              m25_axi_rvalid ,
   output logic                              m25_axi_rready ,
   input  logic [C_M05_AXI_DATA_WIDTH-1:0]   m25_axi_rdata  ,
   input  logic                              m25_axi_rlast  ,

   output logic                              m26_axi_awvalid,
   input  logic                              m26_axi_awready,
   output logic [C_M06_AXI_ADDR_WIDTH-1:0]   m26_axi_awaddr ,
   output logic [8-1:0]                      m26_axi_awlen  ,
   output logic                              m26_axi_wvalid ,
   input  logic                              m26_axi_wready ,
   output logic [C_M06_AXI_DATA_WIDTH-1:0]   m26_axi_wdata  ,
   output logic [C_M06_AXI_DATA_WIDTH/8-1:0] m26_axi_wstrb  ,
   output logic                              m26_axi_wlast  ,
   input  logic                              m26_axi_bvalid ,
   output logic                              m26_axi_bready ,
   output logic                              m26_axi_arvalid,
   input  logic                              m26_axi_arready,
   output logic [C_M06_AXI_ADDR_WIDTH-1:0]   m26_axi_araddr ,
   output logic [8-1:0]                      m26_axi_arlen  ,
   input  logic                              m26_axi_rvalid ,
   output logic                              m26_axi_rready ,
   input  logic [C_M06_AXI_DATA_WIDTH-1:0]   m26_axi_rdata  ,
   input  logic                              m26_axi_rlast  ,

   output logic                              m27_axi_awvalid,
   input  logic                              m27_axi_awready,
   output logic [C_M07_AXI_ADDR_WIDTH-1:0]   m27_axi_awaddr ,
   output logic [8-1:0]                      m27_axi_awlen  ,
   output logic                              m27_axi_wvalid ,
   input  logic                              m27_axi_wready ,
   output logic [C_M07_AXI_DATA_WIDTH-1:0]   m27_axi_wdata  ,
   output logic [C_M07_AXI_DATA_WIDTH/8-1:0] m27_axi_wstrb  ,
   output logic                              m27_axi_wlast  ,
   input  logic                              m27_axi_bvalid ,
   output logic                              m27_axi_bready ,
   output logic                              m27_axi_arvalid,
   input  logic                              m27_axi_arready,
   output logic [C_M07_AXI_ADDR_WIDTH-1:0]   m27_axi_araddr ,
   output logic [8-1:0]                      m27_axi_arlen  ,
   input  logic                              m27_axi_rvalid ,
   output logic                              m27_axi_rready ,
   input  logic [C_M07_AXI_DATA_WIDTH-1:0]   m27_axi_rdata  ,
   input  logic                              m27_axi_rlast  ,

   output logic                              m28_axi_awvalid,
   input  logic                              m28_axi_awready,
   output logic [C_M08_AXI_ADDR_WIDTH-1:0]   m28_axi_awaddr ,
   output logic [8-1:0]                      m28_axi_awlen  ,
   output logic                              m28_axi_wvalid ,
   input  logic                              m28_axi_wready ,
   output logic [C_M08_AXI_DATA_WIDTH-1:0]   m28_axi_wdata  ,
   output logic [C_M08_AXI_DATA_WIDTH/8-1:0] m28_axi_wstrb  ,
   output logic                              m28_axi_wlast  ,
   input  logic                              m28_axi_bvalid ,
   output logic                              m28_axi_bready ,
   output logic                              m28_axi_arvalid,
   input  logic                              m28_axi_arready,
   output logic [C_M08_AXI_ADDR_WIDTH-1:0]   m28_axi_araddr ,
   output logic [8-1:0]                      m28_axi_arlen  ,
   input  logic                              m28_axi_rvalid ,
   output logic                              m28_axi_rready ,
   input  logic [C_M08_AXI_DATA_WIDTH-1:0]   m28_axi_rdata  ,
   input  logic                              m28_axi_rlast  ,

   output logic                              m29_axi_awvalid,
   input  logic                              m29_axi_awready,
   output logic [C_M09_AXI_ADDR_WIDTH-1:0]   m29_axi_awaddr ,
   output logic [8-1:0]                      m29_axi_awlen  ,
   output logic                              m29_axi_wvalid ,
   input  logic                              m29_axi_wready ,
   output logic [C_M09_AXI_DATA_WIDTH-1:0]   m29_axi_wdata  ,
   output logic [C_M09_AXI_DATA_WIDTH/8-1:0] m29_axi_wstrb  ,
   output logic                              m29_axi_wlast  ,
   input  logic                              m29_axi_bvalid ,
   output logic                              m29_axi_bready ,
   output logic                              m29_axi_arvalid,
   input  logic                              m29_axi_arready,
   output logic [C_M09_AXI_ADDR_WIDTH-1:0]   m29_axi_araddr ,
   output logic [8-1:0]                      m29_axi_arlen  ,
   input  logic                              m29_axi_rvalid ,
   output logic                              m29_axi_rready ,
   input  logic [C_M09_AXI_DATA_WIDTH-1:0]   m29_axi_rdata  ,
   input  logic                              m29_axi_rlast  ,

   output logic                              m30_axi_awvalid,
   input  logic                              m30_axi_awready,
   output logic [C_M10_AXI_ADDR_WIDTH-1:0]   m30_axi_awaddr ,
   output logic [8-1:0]                      m30_axi_awlen  ,
   output logic                              m30_axi_wvalid ,
   input  logic                              m30_axi_wready ,
   output logic [C_M10_AXI_DATA_WIDTH-1:0]   m30_axi_wdata  ,
   output logic [C_M10_AXI_DATA_WIDTH/8-1:0] m30_axi_wstrb  ,
   output logic                              m30_axi_wlast  ,
   input  logic                              m30_axi_bvalid ,
   output logic                              m30_axi_bready ,
   output logic                              m30_axi_arvalid,
   input  logic                              m30_axi_arready,
   output logic [C_M10_AXI_ADDR_WIDTH-1:0]   m30_axi_araddr ,
   output logic [8-1:0]                      m30_axi_arlen  ,
   input  logic                              m30_axi_rvalid ,
   output logic                              m30_axi_rready ,
   input  logic [C_M10_AXI_DATA_WIDTH-1:0]   m30_axi_rdata  ,
   input  logic                              m30_axi_rlast  ,

   output logic                              m31_axi_awvalid,
   input  logic                              m31_axi_awready,
   output logic [C_M11_AXI_ADDR_WIDTH-1:0]   m31_axi_awaddr ,
   output logic [8-1:0]                      m31_axi_awlen  ,
   output logic                              m31_axi_wvalid ,
   input  logic                              m31_axi_wready ,
   output logic [C_M11_AXI_DATA_WIDTH-1:0]   m31_axi_wdata  ,
   output logic [C_M11_AXI_DATA_WIDTH/8-1:0] m31_axi_wstrb  ,
   output logic                              m31_axi_wlast  ,
   input  logic                              m31_axi_bvalid ,
   output logic                              m31_axi_bready ,
   output logic                              m31_axi_arvalid,
   input  logic                              m31_axi_arready,
   output logic [C_M11_AXI_ADDR_WIDTH-1:0]   m31_axi_araddr ,
   output logic [8-1:0]                      m31_axi_arlen  ,
   input  logic                              m31_axi_rvalid ,
   output logic                              m31_axi_rready ,
   input  logic [C_M11_AXI_DATA_WIDTH-1:0]   m31_axi_rdata  ,
   input  logic                              m31_axi_rlast  ,

   input  logic [64-1:0]                     axi00_ptr0     ,
   input  logic [64-1:0]                     axi01_ptr0     ,
   input  logic [64-1:0]                     axi02_ptr0     ,
   input  logic [64-1:0]                     axi03_ptr0     ,
   input  logic [64-1:0]                     axi04_ptr0     ,
   input  logic [64-1:0]                     axi05_ptr0     ,
   input  logic [64-1:0]                     axi06_ptr0     ,
   input  logic [64-1:0]                     axi07_ptr0     ,
   input  logic [64-1:0]                     axi08_ptr0     ,
   input  logic [64-1:0]                     axi09_ptr0     ,
   input  logic [64-1:0]                     axi10_ptr0     ,
   input  logic [64-1:0]                     axi11_ptr0     ,
   input  logic [64-1:0]                     axi12_ptr0     ,
   input  logic [64-1:0]                     axi13_ptr0     ,
   input  logic [64-1:0]                     axi14_ptr0     ,
   input  logic [64-1:0]                     axi15_ptr0     ,
   input  logic [64-1:0]                     axi16_ptr0     ,
   input  logic [64-1:0]                     axi17_ptr0     ,
   input  logic [64-1:0]                     axi18_ptr0     ,
   input  logic [64-1:0]                     axi19_ptr0     ,
   input  logic [64-1:0]                     axi20_ptr0     ,
   input  logic [64-1:0]                     axi21_ptr0     ,
   input  logic [64-1:0]                     axi22_ptr0     ,
   input  logic [64-1:0]                     axi23_ptr0     ,
   input  logic [64-1:0]                     axi24_ptr0     ,
   input  logic [64-1:0]                     axi25_ptr0     ,
   input  logic [64-1:0]                     axi26_ptr0     ,
   input  logic [64-1:0]                     axi27_ptr0     ,
   input  logic [64-1:0]                     axi28_ptr0     ,
   input  logic [64-1:0]                     axi29_ptr0     ,
   input  logic [64-1:0]                     axi30_ptr0     ,
   input  logic [64-1:0]                     axi31_ptr0
   );

  logic [2*NLANE-1:0] local_start;
  logic [2*NLANE-1:0] local_done;
  logic [2*NLANE-1:0] local_hold;
  logic [2*NLANE-1:0] local_release;

  always_comb begin
    dbg_ch0_rbeat = '0;
    dbg_ch0_wbeat = '0;
    dbg_ch8_rbeat = '0;
    dbg_ch8_wbeat = '0;
  end

  always_ff @(posedge clk_i) begin
    local_start   <= {NLANE*2{start_i}};
    local_release <= {NLANE*2{local_hold == '1}};
    done_o        <= local_done == '1;
  end

  point_dma_r_channel
    #(
      .ID(0),
      .C_M_AXI_ADDR_WIDTH ( C_M00_AXI_ADDR_WIDTH ),
      .C_M_AXI_DATA_WIDTH ( C_M00_AXI_DATA_WIDTH )
      ) _channel0
      (
       .clk_i,
       .rst_ni,
       .start_i                 ( local_start[0]          ),
       .done_o                  ( local_done[0]           ),
       .hold_o                  ( local_hold[0]           ),
       .release_i               ( local_release[0]        ),
       .we_o                    ( we_o[0]                 ),
       .wdata_o                 ( wdata_o[0]              ),
       .waddr_o                 ( waddr_o[0]              ),
       .wcoarse_o               ( wcoarse_o[0]            ),
       .rcoarse_i               ( rcoarse_i[0]            ),
       .m0_axi_arvalid          ( m00_axi_arvalid         ),
       .m0_axi_arready          ( m00_axi_arready         ),
       .m0_axi_araddr           ( m00_axi_araddr          ),
       .m0_axi_arlen            ( m00_axi_arlen           ),
       .m0_axi_rvalid           ( m00_axi_rvalid          ),
       .m0_axi_rready           ( m00_axi_rready          ),
       .m0_axi_rdata            ( m00_axi_rdata           ),
       .m0_axi_rlast            ( m00_axi_rlast           ),
       .m1_axi_arvalid          ( m01_axi_arvalid         ),
       .m1_axi_arready          ( m01_axi_arready         ),
       .m1_axi_araddr           ( m01_axi_araddr          ),
       .m1_axi_arlen            ( m01_axi_arlen           ),
       .m1_axi_rvalid           ( m01_axi_rvalid          ),
       .m1_axi_rready           ( m01_axi_rready          ),
       .m1_axi_rdata            ( m01_axi_rdata           ),
       .m1_axi_rlast            ( m01_axi_rlast           ),
       .ctrl_addr_offset0       ( axi00_ptr0              ),
       .ctrl_addr_offset1       ( axi01_ptr0              ),
       .dbg_rbeat               (                         ),
       .dbg_rstep               ( dbg_rstep[0]            )
       );

  point_dma_w_channel
    #(
      .ID(1),
      .C_M_AXI_ADDR_WIDTH ( C_M01_AXI_ADDR_WIDTH ),
      .C_M_AXI_DATA_WIDTH ( C_M01_AXI_DATA_WIDTH )
      ) _channel1
      (
       .clk_i,
       .rst_ni,
       .start_i                 ( local_start[1]          ),
       .done_o                  ( local_done[1]           ),
       .hold_o                  ( local_hold[1]           ),
       .release_i               ( local_release[1]        ),
       .re_o                    ( re_o[0]                 ),
       .rdata_i                 ( rdata_i[0]              ),
       .raddr_o                 ( raddr_o[0]              ),
       .wcoarse_i               ( wcoarse_i[0]            ),
       .rcoarse_o               ( rcoarse_o[0]            ),
       .m0_axi_awvalid          ( m00_axi_awvalid         ),
       .m0_axi_awready          ( m00_axi_awready         ),
       .m0_axi_awaddr           ( m00_axi_awaddr          ),
       .m0_axi_awlen            ( m00_axi_awlen           ),
       .m0_axi_wvalid           ( m00_axi_wvalid          ),
       .m0_axi_wready           ( m00_axi_wready          ),
       .m0_axi_wdata            ( m00_axi_wdata           ),
       .m0_axi_wstrb            ( m00_axi_wstrb           ),
       .m0_axi_wlast            ( m00_axi_wlast           ),
       .m0_axi_bvalid           ( m00_axi_bvalid          ),
       .m0_axi_bready           ( m00_axi_bready          ),
       .m1_axi_awvalid          ( m01_axi_awvalid         ),
       .m1_axi_awready          ( m01_axi_awready         ),
       .m1_axi_awaddr           ( m01_axi_awaddr          ),
       .m1_axi_awlen            ( m01_axi_awlen           ),
       .m1_axi_wvalid           ( m01_axi_wvalid          ),
       .m1_axi_wready           ( m01_axi_wready          ),
       .m1_axi_wdata            ( m01_axi_wdata           ),
       .m1_axi_wstrb            ( m01_axi_wstrb           ),
       .m1_axi_wlast            ( m01_axi_wlast           ),
       .m1_axi_bvalid           ( m01_axi_bvalid          ),
       .m1_axi_bready           ( m01_axi_bready          ),
       .ctrl_addr_offset0       ( axi00_ptr0              ),
       .ctrl_addr_offset1       ( axi01_ptr0              ),
       .dbg_wbeat               (                         ),
       .dbg_wstep               ( dbg_wstep[0]            )
       );

  point_dma_r_channel
    #(
      .ID(2),
      .C_M_AXI_ADDR_WIDTH ( C_M02_AXI_ADDR_WIDTH ),
      .C_M_AXI_DATA_WIDTH ( C_M02_AXI_DATA_WIDTH )
      ) _channel2
      (
       .clk_i,
       .rst_ni,
       .start_i                 ( local_start[2]          ),
       .done_o                  ( local_done[2]           ),
       .hold_o                  ( local_hold[2]           ),
       .release_i               ( local_release[2]        ),
       .we_o                    ( we_o[1]                 ),
       .wdata_o                 ( wdata_o[1]              ),
       .waddr_o                 ( waddr_o[1]              ),
       .wcoarse_o               ( wcoarse_o[1]            ),
       .rcoarse_i               ( rcoarse_i[1]            ),
       .m0_axi_arvalid          ( m02_axi_arvalid         ),
       .m0_axi_arready          ( m02_axi_arready         ),
       .m0_axi_araddr           ( m02_axi_araddr          ),
       .m0_axi_arlen            ( m02_axi_arlen           ),
       .m0_axi_rvalid           ( m02_axi_rvalid          ),
       .m0_axi_rready           ( m02_axi_rready          ),
       .m0_axi_rdata            ( m02_axi_rdata           ),
       .m0_axi_rlast            ( m02_axi_rlast           ),
       .m1_axi_arvalid          ( m03_axi_arvalid         ),
       .m1_axi_arready          ( m03_axi_arready         ),
       .m1_axi_araddr           ( m03_axi_araddr          ),
       .m1_axi_arlen            ( m03_axi_arlen           ),
       .m1_axi_rvalid           ( m03_axi_rvalid          ),
       .m1_axi_rready           ( m03_axi_rready          ),
       .m1_axi_rdata            ( m03_axi_rdata           ),
       .m1_axi_rlast            ( m03_axi_rlast           ),
       .ctrl_addr_offset0       ( axi02_ptr0              ),
       .ctrl_addr_offset1       ( axi03_ptr0              ),
       .dbg_rbeat               (                         ),
       .dbg_rstep               ( dbg_rstep[1]            )
       );

  point_dma_w_channel
    #(
      .ID(3),
      .C_M_AXI_ADDR_WIDTH ( C_M03_AXI_ADDR_WIDTH ),
      .C_M_AXI_DATA_WIDTH ( C_M03_AXI_DATA_WIDTH )
      ) _channel3
      (
       .clk_i,
       .rst_ni,
       .start_i                 ( local_start[3]          ),
       .done_o                  ( local_done[3]           ),
       .hold_o                  ( local_hold[3]           ),
       .release_i               ( local_release[3]        ),
       .re_o                    ( re_o[1]                 ),
       .rdata_i                 ( rdata_i[1]              ),
       .raddr_o                 ( raddr_o[1]              ),
       .wcoarse_i               ( wcoarse_i[1]            ),
       .rcoarse_o               ( rcoarse_o[1]            ),
       .m0_axi_awvalid          ( m02_axi_awvalid         ),
       .m0_axi_awready          ( m02_axi_awready         ),
       .m0_axi_awaddr           ( m02_axi_awaddr          ),
       .m0_axi_awlen            ( m02_axi_awlen           ),
       .m0_axi_wvalid           ( m02_axi_wvalid          ),
       .m0_axi_wready           ( m02_axi_wready          ),
       .m0_axi_wdata            ( m02_axi_wdata           ),
       .m0_axi_wstrb            ( m02_axi_wstrb           ),
       .m0_axi_wlast            ( m02_axi_wlast           ),
       .m0_axi_bvalid           ( m02_axi_bvalid          ),
       .m0_axi_bready           ( m02_axi_bready          ),
       .m1_axi_awvalid          ( m03_axi_awvalid         ),
       .m1_axi_awready          ( m03_axi_awready         ),
       .m1_axi_awaddr           ( m03_axi_awaddr          ),
       .m1_axi_awlen            ( m03_axi_awlen           ),
       .m1_axi_wvalid           ( m03_axi_wvalid          ),
       .m1_axi_wready           ( m03_axi_wready          ),
       .m1_axi_wdata            ( m03_axi_wdata           ),
       .m1_axi_wstrb            ( m03_axi_wstrb           ),
       .m1_axi_wlast            ( m03_axi_wlast           ),
       .m1_axi_bvalid           ( m03_axi_bvalid          ),
       .m1_axi_bready           ( m03_axi_bready          ),
       .ctrl_addr_offset0       ( axi02_ptr0              ),
       .ctrl_addr_offset1       ( axi03_ptr0              ),
       .dbg_wbeat               (                         ),
       .dbg_wstep               ( dbg_wstep[1]            )
       );

  point_dma_r_channel
    #(
      .ID(4),
      .C_M_AXI_ADDR_WIDTH ( C_M04_AXI_ADDR_WIDTH ),
      .C_M_AXI_DATA_WIDTH ( C_M04_AXI_DATA_WIDTH )
      ) _channel4
      (
       .clk_i,
       .rst_ni,
       .start_i                 ( local_start[4]          ),
       .done_o                  ( local_done[4]           ),
       .hold_o                  ( local_hold[4]           ),
       .release_i               ( local_release[4]        ),
       .we_o                    ( we_o[2]                 ),
       .wdata_o                 ( wdata_o[2]              ),
       .waddr_o                 ( waddr_o[2]              ),
       .wcoarse_o               ( wcoarse_o[2]            ),
       .rcoarse_i               ( rcoarse_i[2]            ),
       .m0_axi_arvalid          ( m04_axi_arvalid         ),
       .m0_axi_arready          ( m04_axi_arready         ),
       .m0_axi_araddr           ( m04_axi_araddr          ),
       .m0_axi_arlen            ( m04_axi_arlen           ),
       .m0_axi_rvalid           ( m04_axi_rvalid          ),
       .m0_axi_rready           ( m04_axi_rready          ),
       .m0_axi_rdata            ( m04_axi_rdata           ),
       .m0_axi_rlast            ( m04_axi_rlast           ),
       .m1_axi_arvalid          ( m05_axi_arvalid         ),
       .m1_axi_arready          ( m05_axi_arready         ),
       .m1_axi_araddr           ( m05_axi_araddr          ),
       .m1_axi_arlen            ( m05_axi_arlen           ),
       .m1_axi_rvalid           ( m05_axi_rvalid          ),
       .m1_axi_rready           ( m05_axi_rready          ),
       .m1_axi_rdata            ( m05_axi_rdata           ),
       .m1_axi_rlast            ( m05_axi_rlast           ),
       .ctrl_addr_offset0       ( axi04_ptr0              ),
       .ctrl_addr_offset1       ( axi05_ptr0              ),
       .dbg_rbeat               (                         ),
       .dbg_rstep               ( dbg_rstep[2]            )
       );

  point_dma_w_channel
    #(
      .ID(5),
      .C_M_AXI_ADDR_WIDTH ( C_M05_AXI_ADDR_WIDTH ),
      .C_M_AXI_DATA_WIDTH ( C_M05_AXI_DATA_WIDTH )
      ) _channel5
      (
       .clk_i,
       .rst_ni,
       .start_i                 ( local_start[5]          ),
       .done_o                  ( local_done[5]           ),
       .hold_o                  ( local_hold[5]           ),
       .release_i               ( local_release[5]        ),
       .re_o                    ( re_o[2]                 ),
       .rdata_i                 ( rdata_i[2]              ),
       .raddr_o                 ( raddr_o[2]              ),
       .wcoarse_i               ( wcoarse_i[2]            ),
       .rcoarse_o               ( rcoarse_o[2]            ),
       .m0_axi_awvalid          ( m04_axi_awvalid         ),
       .m0_axi_awready          ( m04_axi_awready         ),
       .m0_axi_awaddr           ( m04_axi_awaddr          ),
       .m0_axi_awlen            ( m04_axi_awlen           ),
       .m0_axi_wvalid           ( m04_axi_wvalid          ),
       .m0_axi_wready           ( m04_axi_wready          ),
       .m0_axi_wdata            ( m04_axi_wdata           ),
       .m0_axi_wstrb            ( m04_axi_wstrb           ),
       .m0_axi_wlast            ( m04_axi_wlast           ),
       .m0_axi_bvalid           ( m04_axi_bvalid          ),
       .m0_axi_bready           ( m04_axi_bready          ),
       .m1_axi_awvalid          ( m05_axi_awvalid         ),
       .m1_axi_awready          ( m05_axi_awready         ),
       .m1_axi_awaddr           ( m05_axi_awaddr          ),
       .m1_axi_awlen            ( m05_axi_awlen           ),
       .m1_axi_wvalid           ( m05_axi_wvalid          ),
       .m1_axi_wready           ( m05_axi_wready          ),
       .m1_axi_wdata            ( m05_axi_wdata           ),
       .m1_axi_wstrb            ( m05_axi_wstrb           ),
       .m1_axi_wlast            ( m05_axi_wlast           ),
       .m1_axi_bvalid           ( m05_axi_bvalid          ),
       .m1_axi_bready           ( m05_axi_bready          ),
       .ctrl_addr_offset0       ( axi04_ptr0              ),
       .ctrl_addr_offset1       ( axi05_ptr0              ),
       .dbg_wbeat               (                         ),
       .dbg_wstep               ( dbg_wstep[2]            )
       );

  point_dma_r_channel
    #(
      .ID(6),
      .C_M_AXI_ADDR_WIDTH ( C_M06_AXI_ADDR_WIDTH ),
      .C_M_AXI_DATA_WIDTH ( C_M06_AXI_DATA_WIDTH )
      ) _channel6
      (
       .clk_i,
       .rst_ni,
       .start_i                 ( local_start[6]          ),
       .done_o                  ( local_done[6]           ),
       .hold_o                  ( local_hold[6]           ),
       .release_i               ( local_release[6]        ),
       .we_o                    ( we_o[3]                 ),
       .wdata_o                 ( wdata_o[3]              ),
       .waddr_o                 ( waddr_o[3]              ),
       .wcoarse_o               ( wcoarse_o[3]            ),
       .rcoarse_i               ( rcoarse_i[3]            ),
       .m0_axi_arvalid          ( m06_axi_arvalid         ),
       .m0_axi_arready          ( m06_axi_arready         ),
       .m0_axi_araddr           ( m06_axi_araddr          ),
       .m0_axi_arlen            ( m06_axi_arlen           ),
       .m0_axi_rvalid           ( m06_axi_rvalid          ),
       .m0_axi_rready           ( m06_axi_rready          ),
       .m0_axi_rdata            ( m06_axi_rdata           ),
       .m0_axi_rlast            ( m06_axi_rlast           ),
       .m1_axi_arvalid          ( m07_axi_arvalid         ),
       .m1_axi_arready          ( m07_axi_arready         ),
       .m1_axi_araddr           ( m07_axi_araddr          ),
       .m1_axi_arlen            ( m07_axi_arlen           ),
       .m1_axi_rvalid           ( m07_axi_rvalid          ),
       .m1_axi_rready           ( m07_axi_rready          ),
       .m1_axi_rdata            ( m07_axi_rdata           ),
       .m1_axi_rlast            ( m07_axi_rlast           ),
       .ctrl_addr_offset0       ( axi06_ptr0              ),
       .ctrl_addr_offset1       ( axi07_ptr0              ),
       .dbg_rbeat               (                         ),
       .dbg_rstep               ( dbg_rstep[3]            )
       );

  point_dma_w_channel
    #(
      .ID(7),
      .C_M_AXI_ADDR_WIDTH ( C_M07_AXI_ADDR_WIDTH ),
      .C_M_AXI_DATA_WIDTH ( C_M07_AXI_DATA_WIDTH )
      ) _channel7
      (
       .clk_i,
       .rst_ni,
       .start_i                 ( local_start[7]          ),
       .done_o                  ( local_done[7]           ),
       .hold_o                  ( local_hold[7]           ),
       .release_i               ( local_release[7]        ),
       .re_o                    ( re_o[3]                 ),
       .rdata_i                 ( rdata_i[3]              ),
       .raddr_o                 ( raddr_o[3]              ),
       .wcoarse_i               ( wcoarse_i[3]            ),
       .rcoarse_o               ( rcoarse_o[3]            ),
       .m0_axi_awvalid          ( m06_axi_awvalid         ),
       .m0_axi_awready          ( m06_axi_awready         ),
       .m0_axi_awaddr           ( m06_axi_awaddr          ),
       .m0_axi_awlen            ( m06_axi_awlen           ),
       .m0_axi_wvalid           ( m06_axi_wvalid          ),
       .m0_axi_wready           ( m06_axi_wready          ),
       .m0_axi_wdata            ( m06_axi_wdata           ),
       .m0_axi_wstrb            ( m06_axi_wstrb           ),
       .m0_axi_wlast            ( m06_axi_wlast           ),
       .m0_axi_bvalid           ( m06_axi_bvalid          ),
       .m0_axi_bready           ( m06_axi_bready          ),
       .m1_axi_awvalid          ( m07_axi_awvalid         ),
       .m1_axi_awready          ( m07_axi_awready         ),
       .m1_axi_awaddr           ( m07_axi_awaddr          ),
       .m1_axi_awlen            ( m07_axi_awlen           ),
       .m1_axi_wvalid           ( m07_axi_wvalid          ),
       .m1_axi_wready           ( m07_axi_wready          ),
       .m1_axi_wdata            ( m07_axi_wdata           ),
       .m1_axi_wstrb            ( m07_axi_wstrb           ),
       .m1_axi_wlast            ( m07_axi_wlast           ),
       .m1_axi_bvalid           ( m07_axi_bvalid          ),
       .m1_axi_bready           ( m07_axi_bready          ),
       .ctrl_addr_offset0       ( axi06_ptr0              ),
       .ctrl_addr_offset1       ( axi07_ptr0              ),
       .dbg_wbeat               (                         ),
       .dbg_wstep               ( dbg_wstep[3]            )
       );

  point_dma_r_channel
    #(
      .ID(8),
      .C_M_AXI_ADDR_WIDTH ( C_M08_AXI_ADDR_WIDTH ),
      .C_M_AXI_DATA_WIDTH ( C_M08_AXI_DATA_WIDTH )
      ) _channel8
      (
       .clk_i,
       .rst_ni,
       .start_i                 ( local_start[8]          ),
       .done_o                  ( local_done[8]           ),
       .hold_o                  ( local_hold[8]           ),
       .release_i               ( local_release[8]        ),
       .we_o                    ( we_o[4]                 ),
       .wdata_o                 ( wdata_o[4]              ),
       .waddr_o                 ( waddr_o[4]              ),
       .wcoarse_o               ( wcoarse_o[4]            ),
       .rcoarse_i               ( rcoarse_i[4]            ),
       .m0_axi_arvalid          ( m08_axi_arvalid         ),
       .m0_axi_arready          ( m08_axi_arready         ),
       .m0_axi_araddr           ( m08_axi_araddr          ),
       .m0_axi_arlen            ( m08_axi_arlen           ),
       .m0_axi_rvalid           ( m08_axi_rvalid          ),
       .m0_axi_rready           ( m08_axi_rready          ),
       .m0_axi_rdata            ( m08_axi_rdata           ),
       .m0_axi_rlast            ( m08_axi_rlast           ),
       .m1_axi_arvalid          ( m09_axi_arvalid         ),
       .m1_axi_arready          ( m09_axi_arready         ),
       .m1_axi_araddr           ( m09_axi_araddr          ),
       .m1_axi_arlen            ( m09_axi_arlen           ),
       .m1_axi_rvalid           ( m09_axi_rvalid          ),
       .m1_axi_rready           ( m09_axi_rready          ),
       .m1_axi_rdata            ( m09_axi_rdata           ),
       .m1_axi_rlast            ( m09_axi_rlast           ),
       .ctrl_addr_offset0       ( axi08_ptr0              ),
       .ctrl_addr_offset1       ( axi09_ptr0              ),
       .dbg_rbeat               (                         ),
       .dbg_rstep               ( dbg_rstep[4]            )
       );

  point_dma_w_channel
    #(
      .ID(9),
      .C_M_AXI_ADDR_WIDTH ( C_M09_AXI_ADDR_WIDTH ),
      .C_M_AXI_DATA_WIDTH ( C_M09_AXI_DATA_WIDTH )
      ) _channel9
      (
       .clk_i,
       .rst_ni,
       .start_i                 ( local_start[9]          ),
       .done_o                  ( local_done[9]           ),
       .hold_o                  ( local_hold[9]           ),
       .release_i               ( local_release[9]        ),
       .re_o                    ( re_o[4]                 ),
       .rdata_i                 ( rdata_i[4]              ),
       .raddr_o                 ( raddr_o[4]              ),
       .wcoarse_i               ( wcoarse_i[4]            ),
       .rcoarse_o               ( rcoarse_o[4]            ),
       .m0_axi_awvalid          ( m08_axi_awvalid         ),
       .m0_axi_awready          ( m08_axi_awready         ),
       .m0_axi_awaddr           ( m08_axi_awaddr          ),
       .m0_axi_awlen            ( m08_axi_awlen           ),
       .m0_axi_wvalid           ( m08_axi_wvalid          ),
       .m0_axi_wready           ( m08_axi_wready          ),
       .m0_axi_wdata            ( m08_axi_wdata           ),
       .m0_axi_wstrb            ( m08_axi_wstrb           ),
       .m0_axi_wlast            ( m08_axi_wlast           ),
       .m0_axi_bvalid           ( m08_axi_bvalid          ),
       .m0_axi_bready           ( m08_axi_bready          ),
       .m1_axi_awvalid          ( m09_axi_awvalid         ),
       .m1_axi_awready          ( m09_axi_awready         ),
       .m1_axi_awaddr           ( m09_axi_awaddr          ),
       .m1_axi_awlen            ( m09_axi_awlen           ),
       .m1_axi_wvalid           ( m09_axi_wvalid          ),
       .m1_axi_wready           ( m09_axi_wready          ),
       .m1_axi_wdata            ( m09_axi_wdata           ),
       .m1_axi_wstrb            ( m09_axi_wstrb           ),
       .m1_axi_wlast            ( m09_axi_wlast           ),
       .m1_axi_bvalid           ( m09_axi_bvalid          ),
       .m1_axi_bready           ( m09_axi_bready          ),
       .ctrl_addr_offset0       ( axi08_ptr0              ),
       .ctrl_addr_offset1       ( axi09_ptr0              ),
       .dbg_wbeat               (                         ),
       .dbg_wstep               ( dbg_wstep[4]            )
       );

  point_dma_r_channel
    #(
      .ID(10),
      .C_M_AXI_ADDR_WIDTH ( C_M10_AXI_ADDR_WIDTH ),
      .C_M_AXI_DATA_WIDTH ( C_M10_AXI_DATA_WIDTH )
      ) _channel10
      (
       .clk_i,
       .rst_ni,
       .start_i                 ( local_start[10]         ),
       .done_o                  ( local_done[10]          ),
       .hold_o                  ( local_hold[10]          ),
       .release_i               ( local_release[10]       ),
       .we_o                    ( we_o[5]                 ),
       .wdata_o                 ( wdata_o[5]              ),
       .waddr_o                 ( waddr_o[5]              ),
       .wcoarse_o               ( wcoarse_o[5]            ),
       .rcoarse_i               ( rcoarse_i[5]            ),
       .m0_axi_arvalid          ( m10_axi_arvalid         ),
       .m0_axi_arready          ( m10_axi_arready         ),
       .m0_axi_araddr           ( m10_axi_araddr          ),
       .m0_axi_arlen            ( m10_axi_arlen           ),
       .m0_axi_rvalid           ( m10_axi_rvalid          ),
       .m0_axi_rready           ( m10_axi_rready          ),
       .m0_axi_rdata            ( m10_axi_rdata           ),
       .m0_axi_rlast            ( m10_axi_rlast           ),
       .m1_axi_arvalid          ( m11_axi_arvalid         ),
       .m1_axi_arready          ( m11_axi_arready         ),
       .m1_axi_araddr           ( m11_axi_araddr          ),
       .m1_axi_arlen            ( m11_axi_arlen           ),
       .m1_axi_rvalid           ( m11_axi_rvalid          ),
       .m1_axi_rready           ( m11_axi_rready          ),
       .m1_axi_rdata            ( m11_axi_rdata           ),
       .m1_axi_rlast            ( m11_axi_rlast           ),
       .ctrl_addr_offset0       ( axi10_ptr0              ),
       .ctrl_addr_offset1       ( axi11_ptr0              ),
       .dbg_rbeat               (                         ),
       .dbg_rstep               ( dbg_rstep[5]            )
       );

  point_dma_w_channel
    #(
      .ID(11),
      .C_M_AXI_ADDR_WIDTH ( C_M11_AXI_ADDR_WIDTH ),
      .C_M_AXI_DATA_WIDTH ( C_M11_AXI_DATA_WIDTH )
      ) _channel11
      (
       .clk_i,
       .rst_ni,
       .start_i                 ( local_start[11]         ),
       .done_o                  ( local_done[11]          ),
       .hold_o                  ( local_hold[11]          ),
       .release_i               ( local_release[11]       ),
       .re_o                    ( re_o[5]                 ),
       .rdata_i                 ( rdata_i[5]              ),
       .raddr_o                 ( raddr_o[5]              ),
       .wcoarse_i               ( wcoarse_i[5]            ),
       .rcoarse_o               ( rcoarse_o[5]            ),
       .m0_axi_awvalid          ( m10_axi_awvalid         ),
       .m0_axi_awready          ( m10_axi_awready         ),
       .m0_axi_awaddr           ( m10_axi_awaddr          ),
       .m0_axi_awlen            ( m10_axi_awlen           ),
       .m0_axi_wvalid           ( m10_axi_wvalid          ),
       .m0_axi_wready           ( m10_axi_wready          ),
       .m0_axi_wdata            ( m10_axi_wdata           ),
       .m0_axi_wstrb            ( m10_axi_wstrb           ),
       .m0_axi_wlast            ( m10_axi_wlast           ),
       .m0_axi_bvalid           ( m10_axi_bvalid          ),
       .m0_axi_bready           ( m10_axi_bready          ),
       .m1_axi_awvalid          ( m11_axi_awvalid         ),
       .m1_axi_awready          ( m11_axi_awready         ),
       .m1_axi_awaddr           ( m11_axi_awaddr          ),
       .m1_axi_awlen            ( m11_axi_awlen           ),
       .m1_axi_wvalid           ( m11_axi_wvalid          ),
       .m1_axi_wready           ( m11_axi_wready          ),
       .m1_axi_wdata            ( m11_axi_wdata           ),
       .m1_axi_wstrb            ( m11_axi_wstrb           ),
       .m1_axi_wlast            ( m11_axi_wlast           ),
       .m1_axi_bvalid           ( m11_axi_bvalid          ),
       .m1_axi_bready           ( m11_axi_bready          ),
       .ctrl_addr_offset0       ( axi10_ptr0              ),
       .ctrl_addr_offset1       ( axi11_ptr0              ),
       .dbg_wbeat               (                         ),
       .dbg_wstep               ( dbg_wstep[5]            )
       );

  point_dma_r_channel
    #(
      .ID(12),
      .C_M_AXI_ADDR_WIDTH ( C_M12_AXI_ADDR_WIDTH ),
      .C_M_AXI_DATA_WIDTH ( C_M12_AXI_DATA_WIDTH )
      ) _channel12
      (
       .clk_i,
       .rst_ni,
       .start_i                 ( local_start[12]         ),
       .done_o                  ( local_done[12]          ),
       .hold_o                  ( local_hold[12]          ),
       .release_i               ( local_release[12]       ),
       .we_o                    ( we_o[6]                 ),
       .wdata_o                 ( wdata_o[6]              ),
       .waddr_o                 ( waddr_o[6]              ),
       .wcoarse_o               ( wcoarse_o[6]            ),
       .rcoarse_i               ( rcoarse_i[6]            ),
       .m0_axi_arvalid          ( m12_axi_arvalid         ),
       .m0_axi_arready          ( m12_axi_arready         ),
       .m0_axi_araddr           ( m12_axi_araddr          ),
       .m0_axi_arlen            ( m12_axi_arlen           ),
       .m0_axi_rvalid           ( m12_axi_rvalid          ),
       .m0_axi_rready           ( m12_axi_rready          ),
       .m0_axi_rdata            ( m12_axi_rdata           ),
       .m0_axi_rlast            ( m12_axi_rlast           ),
       .m1_axi_arvalid          ( m13_axi_arvalid         ),
       .m1_axi_arready          ( m13_axi_arready         ),
       .m1_axi_araddr           ( m13_axi_araddr          ),
       .m1_axi_arlen            ( m13_axi_arlen           ),
       .m1_axi_rvalid           ( m13_axi_rvalid          ),
       .m1_axi_rready           ( m13_axi_rready          ),
       .m1_axi_rdata            ( m13_axi_rdata           ),
       .m1_axi_rlast            ( m13_axi_rlast           ),
       .ctrl_addr_offset0       ( axi12_ptr0              ),
       .ctrl_addr_offset1       ( axi13_ptr0              ),
       .dbg_rbeat               (                         ),
       .dbg_rstep               ( dbg_rstep[6]            )
       );

  point_dma_w_channel
    #(
      .ID(13),
      .C_M_AXI_ADDR_WIDTH ( C_M13_AXI_ADDR_WIDTH ),
      .C_M_AXI_DATA_WIDTH ( C_M13_AXI_DATA_WIDTH )
      ) _channel13
      (
       .clk_i,
       .rst_ni,
       .start_i                 ( local_start[13]         ),
       .done_o                  ( local_done[13]          ),
       .hold_o                  ( local_hold[13]          ),
       .release_i               ( local_release[13]       ),
       .re_o                    ( re_o[6]                 ),
       .rdata_i                 ( rdata_i[6]              ),
       .raddr_o                 ( raddr_o[6]              ),
       .wcoarse_i               ( wcoarse_i[6]            ),
       .rcoarse_o               ( rcoarse_o[6]            ),
       .m0_axi_awvalid          ( m12_axi_awvalid         ),
       .m0_axi_awready          ( m12_axi_awready         ),
       .m0_axi_awaddr           ( m12_axi_awaddr          ),
       .m0_axi_awlen            ( m12_axi_awlen           ),
       .m0_axi_wvalid           ( m12_axi_wvalid          ),
       .m0_axi_wready           ( m12_axi_wready          ),
       .m0_axi_wdata            ( m12_axi_wdata           ),
       .m0_axi_wstrb            ( m12_axi_wstrb           ),
       .m0_axi_wlast            ( m12_axi_wlast           ),
       .m0_axi_bvalid           ( m12_axi_bvalid          ),
       .m0_axi_bready           ( m12_axi_bready          ),
       .m1_axi_awvalid          ( m13_axi_awvalid         ),
       .m1_axi_awready          ( m13_axi_awready         ),
       .m1_axi_awaddr           ( m13_axi_awaddr          ),
       .m1_axi_awlen            ( m13_axi_awlen           ),
       .m1_axi_wvalid           ( m13_axi_wvalid          ),
       .m1_axi_wready           ( m13_axi_wready          ),
       .m1_axi_wdata            ( m13_axi_wdata           ),
       .m1_axi_wstrb            ( m13_axi_wstrb           ),
       .m1_axi_wlast            ( m13_axi_wlast           ),
       .m1_axi_bvalid           ( m13_axi_bvalid          ),
       .m1_axi_bready           ( m13_axi_bready          ),
       .ctrl_addr_offset0       ( axi12_ptr0              ),
       .ctrl_addr_offset1       ( axi13_ptr0              ),
       .dbg_wbeat               (                         ),
       .dbg_wstep               ( dbg_wstep[6]            )
       );

  point_dma_r_channel
    #(
      .ID(14),
      .C_M_AXI_ADDR_WIDTH ( C_M14_AXI_ADDR_WIDTH ),
      .C_M_AXI_DATA_WIDTH ( C_M14_AXI_DATA_WIDTH )
      ) _channel14
      (
       .clk_i,
       .rst_ni,
       .start_i                 ( local_start[14]         ),
       .done_o                  ( local_done[14]          ),
       .hold_o                  ( local_hold[14]          ),
       .release_i               ( local_release[14]       ),
       .we_o                    ( we_o[7]                 ),
       .wdata_o                 ( wdata_o[7]              ),
       .waddr_o                 ( waddr_o[7]              ),
       .wcoarse_o               ( wcoarse_o[7]            ),
       .rcoarse_i               ( rcoarse_i[7]            ),
       .m0_axi_arvalid          ( m14_axi_arvalid         ),
       .m0_axi_arready          ( m14_axi_arready         ),
       .m0_axi_araddr           ( m14_axi_araddr          ),
       .m0_axi_arlen            ( m14_axi_arlen           ),
       .m0_axi_rvalid           ( m14_axi_rvalid          ),
       .m0_axi_rready           ( m14_axi_rready          ),
       .m0_axi_rdata            ( m14_axi_rdata           ),
       .m0_axi_rlast            ( m14_axi_rlast           ),
       .m1_axi_arvalid          ( m15_axi_arvalid         ),
       .m1_axi_arready          ( m15_axi_arready         ),
       .m1_axi_araddr           ( m15_axi_araddr          ),
       .m1_axi_arlen            ( m15_axi_arlen           ),
       .m1_axi_rvalid           ( m15_axi_rvalid          ),
       .m1_axi_rready           ( m15_axi_rready          ),
       .m1_axi_rdata            ( m15_axi_rdata           ),
       .m1_axi_rlast            ( m15_axi_rlast           ),
       .ctrl_addr_offset0       ( axi14_ptr0              ),
       .ctrl_addr_offset1       ( axi15_ptr0              ),
       .dbg_rbeat               (                         ),
       .dbg_rstep               ( dbg_rstep[7]            )
       );

  point_dma_w_channel
    #(
      .ID(15),
      .C_M_AXI_ADDR_WIDTH ( C_M15_AXI_ADDR_WIDTH ),
      .C_M_AXI_DATA_WIDTH ( C_M15_AXI_DATA_WIDTH )
      ) _channel15
      (
       .clk_i,
       .rst_ni,
       .start_i                 ( local_start[15]         ),
       .done_o                  ( local_done[15]          ),
       .hold_o                  ( local_hold[15]          ),
       .release_i               ( local_release[15]       ),
       .re_o                    ( re_o[7]                 ),
       .rdata_i                 ( rdata_i[7]              ),
       .raddr_o                 ( raddr_o[7]              ),
       .wcoarse_i               ( wcoarse_i[7]            ),
       .rcoarse_o               ( rcoarse_o[7]            ),
       .m0_axi_awvalid          ( m14_axi_awvalid         ),
       .m0_axi_awready          ( m14_axi_awready         ),
       .m0_axi_awaddr           ( m14_axi_awaddr          ),
       .m0_axi_awlen            ( m14_axi_awlen           ),
       .m0_axi_wvalid           ( m14_axi_wvalid          ),
       .m0_axi_wready           ( m14_axi_wready          ),
       .m0_axi_wdata            ( m14_axi_wdata           ),
       .m0_axi_wstrb            ( m14_axi_wstrb           ),
       .m0_axi_wlast            ( m14_axi_wlast           ),
       .m0_axi_bvalid           ( m14_axi_bvalid          ),
       .m0_axi_bready           ( m14_axi_bready          ),
       .m1_axi_awvalid          ( m15_axi_awvalid         ),
       .m1_axi_awready          ( m15_axi_awready         ),
       .m1_axi_awaddr           ( m15_axi_awaddr          ),
       .m1_axi_awlen            ( m15_axi_awlen           ),
       .m1_axi_wvalid           ( m15_axi_wvalid          ),
       .m1_axi_wready           ( m15_axi_wready          ),
       .m1_axi_wdata            ( m15_axi_wdata           ),
       .m1_axi_wstrb            ( m15_axi_wstrb           ),
       .m1_axi_wlast            ( m15_axi_wlast           ),
       .m1_axi_bvalid           ( m15_axi_bvalid          ),
       .m1_axi_bready           ( m15_axi_bready          ),
       .ctrl_addr_offset0       ( axi14_ptr0              ),
       .ctrl_addr_offset1       ( axi15_ptr0              ),
       .dbg_wbeat               (                         ),
       .dbg_wstep               ( dbg_wstep[7]            )
       );

  point_dma_r_channel
    #(
      .ID(16),
      .C_M_AXI_ADDR_WIDTH ( C_M16_AXI_ADDR_WIDTH ),
      .C_M_AXI_DATA_WIDTH ( C_M16_AXI_DATA_WIDTH )
      ) _channel16
      (
       .clk_i,
       .rst_ni,
       .start_i                 ( local_start[16]         ),
       .done_o                  ( local_done[16]          ),
       .hold_o                  ( local_hold[16]          ),
       .release_i               ( local_release[16]       ),
       .we_o                    ( we_o[8]                 ),
       .wdata_o                 ( wdata_o[8]              ),
       .waddr_o                 ( waddr_o[8]              ),
       .wcoarse_o               ( wcoarse_o[8]            ),
       .rcoarse_i               ( rcoarse_i[8]            ),
       .m0_axi_arvalid          ( m16_axi_arvalid         ),
       .m0_axi_arready          ( m16_axi_arready         ),
       .m0_axi_araddr           ( m16_axi_araddr          ),
       .m0_axi_arlen            ( m16_axi_arlen           ),
       .m0_axi_rvalid           ( m16_axi_rvalid          ),
       .m0_axi_rready           ( m16_axi_rready          ),
       .m0_axi_rdata            ( m16_axi_rdata           ),
       .m0_axi_rlast            ( m16_axi_rlast           ),
       .m1_axi_arvalid          ( m17_axi_arvalid         ),
       .m1_axi_arready          ( m17_axi_arready         ),
       .m1_axi_araddr           ( m17_axi_araddr          ),
       .m1_axi_arlen            ( m17_axi_arlen           ),
       .m1_axi_rvalid           ( m17_axi_rvalid          ),
       .m1_axi_rready           ( m17_axi_rready          ),
       .m1_axi_rdata            ( m17_axi_rdata           ),
       .m1_axi_rlast            ( m17_axi_rlast           ),
       .ctrl_addr_offset0       ( axi16_ptr0              ),
       .ctrl_addr_offset1       ( axi17_ptr0              ),
       .dbg_rbeat               (                         ),
       .dbg_rstep               ( dbg_rstep[8]            )
       );

  point_dma_w_channel
    #(
      .ID(17),
      .C_M_AXI_ADDR_WIDTH ( C_M17_AXI_ADDR_WIDTH ),
      .C_M_AXI_DATA_WIDTH ( C_M17_AXI_DATA_WIDTH )
      ) _channel17
      (
       .clk_i,
       .rst_ni,
       .start_i                 ( local_start[17]         ),
       .done_o                  ( local_done[17]          ),
       .hold_o                  ( local_hold[17]          ),
       .release_i               ( local_release[17]       ),
       .re_o                    ( re_o[8]                 ),
       .rdata_i                 ( rdata_i[8]              ),
       .raddr_o                 ( raddr_o[8]              ),
       .wcoarse_i               ( wcoarse_i[8]            ),
       .rcoarse_o               ( rcoarse_o[8]            ),
       .m0_axi_awvalid          ( m16_axi_awvalid         ),
       .m0_axi_awready          ( m16_axi_awready         ),
       .m0_axi_awaddr           ( m16_axi_awaddr          ),
       .m0_axi_awlen            ( m16_axi_awlen           ),
       .m0_axi_wvalid           ( m16_axi_wvalid          ),
       .m0_axi_wready           ( m16_axi_wready          ),
       .m0_axi_wdata            ( m16_axi_wdata           ),
       .m0_axi_wstrb            ( m16_axi_wstrb           ),
       .m0_axi_wlast            ( m16_axi_wlast           ),
       .m0_axi_bvalid           ( m16_axi_bvalid          ),
       .m0_axi_bready           ( m16_axi_bready          ),
       .m1_axi_awvalid          ( m17_axi_awvalid         ),
       .m1_axi_awready          ( m17_axi_awready         ),
       .m1_axi_awaddr           ( m17_axi_awaddr          ),
       .m1_axi_awlen            ( m17_axi_awlen           ),
       .m1_axi_wvalid           ( m17_axi_wvalid          ),
       .m1_axi_wready           ( m17_axi_wready          ),
       .m1_axi_wdata            ( m17_axi_wdata           ),
       .m1_axi_wstrb            ( m17_axi_wstrb           ),
       .m1_axi_wlast            ( m17_axi_wlast           ),
       .m1_axi_bvalid           ( m17_axi_bvalid          ),
       .m1_axi_bready           ( m17_axi_bready          ),
       .ctrl_addr_offset0       ( axi16_ptr0              ),
       .ctrl_addr_offset1       ( axi17_ptr0              ),
       .dbg_wbeat               (                         ),
       .dbg_wstep               ( dbg_wstep[8]            )
       );

  point_dma_r_channel
    #(
      .ID(18),
      .C_M_AXI_ADDR_WIDTH ( C_M18_AXI_ADDR_WIDTH ),
      .C_M_AXI_DATA_WIDTH ( C_M18_AXI_DATA_WIDTH )
      ) _channel18
      (
       .clk_i,
       .rst_ni,
       .start_i                 ( local_start[18]         ),
       .done_o                  ( local_done[18]          ),
       .hold_o                  ( local_hold[18]          ),
       .release_i               ( local_release[18]       ),
       .we_o                    ( we_o[9]                 ),
       .wdata_o                 ( wdata_o[9]              ),
       .waddr_o                 ( waddr_o[9]              ),
       .wcoarse_o               ( wcoarse_o[9]            ),
       .rcoarse_i               ( rcoarse_i[9]            ),
       .m0_axi_arvalid          ( m18_axi_arvalid         ),
       .m0_axi_arready          ( m18_axi_arready         ),
       .m0_axi_araddr           ( m18_axi_araddr          ),
       .m0_axi_arlen            ( m18_axi_arlen           ),
       .m0_axi_rvalid           ( m18_axi_rvalid          ),
       .m0_axi_rready           ( m18_axi_rready          ),
       .m0_axi_rdata            ( m18_axi_rdata           ),
       .m0_axi_rlast            ( m18_axi_rlast           ),
       .m1_axi_arvalid          ( m19_axi_arvalid         ),
       .m1_axi_arready          ( m19_axi_arready         ),
       .m1_axi_araddr           ( m19_axi_araddr          ),
       .m1_axi_arlen            ( m19_axi_arlen           ),
       .m1_axi_rvalid           ( m19_axi_rvalid          ),
       .m1_axi_rready           ( m19_axi_rready          ),
       .m1_axi_rdata            ( m19_axi_rdata           ),
       .m1_axi_rlast            ( m19_axi_rlast           ),
       .ctrl_addr_offset0       ( axi18_ptr0              ),
       .ctrl_addr_offset1       ( axi19_ptr0              ),
       .dbg_rbeat               (                         ),
       .dbg_rstep               ( dbg_rstep[9]            )
       );

  point_dma_w_channel
    #(
      .ID(19),
      .C_M_AXI_ADDR_WIDTH ( C_M19_AXI_ADDR_WIDTH ),
      .C_M_AXI_DATA_WIDTH ( C_M19_AXI_DATA_WIDTH )
      ) _channel19
      (
       .clk_i,
       .rst_ni,
       .start_i                 ( local_start[19]         ),
       .done_o                  ( local_done[19]          ),
       .hold_o                  ( local_hold[19]          ),
       .release_i               ( local_release[19]       ),
       .re_o                    ( re_o[9]                 ),
       .rdata_i                 ( rdata_i[9]              ),
       .raddr_o                 ( raddr_o[9]              ),
       .wcoarse_i               ( wcoarse_i[9]            ),
       .rcoarse_o               ( rcoarse_o[9]            ),
       .m0_axi_awvalid          ( m18_axi_awvalid         ),
       .m0_axi_awready          ( m18_axi_awready         ),
       .m0_axi_awaddr           ( m18_axi_awaddr          ),
       .m0_axi_awlen            ( m18_axi_awlen           ),
       .m0_axi_wvalid           ( m18_axi_wvalid          ),
       .m0_axi_wready           ( m18_axi_wready          ),
       .m0_axi_wdata            ( m18_axi_wdata           ),
       .m0_axi_wstrb            ( m18_axi_wstrb           ),
       .m0_axi_wlast            ( m18_axi_wlast           ),
       .m0_axi_bvalid           ( m18_axi_bvalid          ),
       .m0_axi_bready           ( m18_axi_bready          ),
       .m1_axi_awvalid          ( m19_axi_awvalid         ),
       .m1_axi_awready          ( m19_axi_awready         ),
       .m1_axi_awaddr           ( m19_axi_awaddr          ),
       .m1_axi_awlen            ( m19_axi_awlen           ),
       .m1_axi_wvalid           ( m19_axi_wvalid          ),
       .m1_axi_wready           ( m19_axi_wready          ),
       .m1_axi_wdata            ( m19_axi_wdata           ),
       .m1_axi_wstrb            ( m19_axi_wstrb           ),
       .m1_axi_wlast            ( m19_axi_wlast           ),
       .m1_axi_bvalid           ( m19_axi_bvalid          ),
       .m1_axi_bready           ( m19_axi_bready          ),
       .ctrl_addr_offset0       ( axi18_ptr0              ),
       .ctrl_addr_offset1       ( axi19_ptr0              ),
       .dbg_wbeat               (                         ),
       .dbg_wstep               ( dbg_wstep[9]            )
       );

  point_dma_r_channel
    #(
      .ID(20),
      .C_M_AXI_ADDR_WIDTH ( C_M20_AXI_ADDR_WIDTH ),
      .C_M_AXI_DATA_WIDTH ( C_M20_AXI_DATA_WIDTH )
      ) _channel20
      (
       .clk_i,
       .rst_ni,
       .start_i                 ( local_start[20]         ),
       .done_o                  ( local_done[20]          ),
       .hold_o                  ( local_hold[20]          ),
       .release_i               ( local_release[20]       ),
       .we_o                    ( we_o[10]                ),
       .wdata_o                 ( wdata_o[10]             ),
       .waddr_o                 ( waddr_o[10]             ),
       .wcoarse_o               ( wcoarse_o[10]           ),
       .rcoarse_i               ( rcoarse_i[10]           ),
       .m0_axi_arvalid          ( m20_axi_arvalid         ),
       .m0_axi_arready          ( m20_axi_arready         ),
       .m0_axi_araddr           ( m20_axi_araddr          ),
       .m0_axi_arlen            ( m20_axi_arlen           ),
       .m0_axi_rvalid           ( m20_axi_rvalid          ),
       .m0_axi_rready           ( m20_axi_rready          ),
       .m0_axi_rdata            ( m20_axi_rdata           ),
       .m0_axi_rlast            ( m20_axi_rlast           ),
       .m1_axi_arvalid          ( m21_axi_arvalid         ),
       .m1_axi_arready          ( m21_axi_arready         ),
       .m1_axi_araddr           ( m21_axi_araddr          ),
       .m1_axi_arlen            ( m21_axi_arlen           ),
       .m1_axi_rvalid           ( m21_axi_rvalid          ),
       .m1_axi_rready           ( m21_axi_rready          ),
       .m1_axi_rdata            ( m21_axi_rdata           ),
       .m1_axi_rlast            ( m21_axi_rlast           ),
       .ctrl_addr_offset0       ( axi20_ptr0              ),
       .ctrl_addr_offset1       ( axi21_ptr0              ),
       .dbg_rbeat               (                         ),
       .dbg_rstep               ( dbg_rstep[10]           )
       );

  point_dma_w_channel
    #(
      .ID(21),
      .C_M_AXI_ADDR_WIDTH ( C_M21_AXI_ADDR_WIDTH ),
      .C_M_AXI_DATA_WIDTH ( C_M21_AXI_DATA_WIDTH )
      ) _channel21
      (
       .clk_i,
       .rst_ni,
       .start_i                 ( local_start[21]         ),
       .done_o                  ( local_done[21]          ),
       .hold_o                  ( local_hold[21]          ),
       .release_i               ( local_release[21]       ),
       .re_o                    ( re_o[10]                ),
       .rdata_i                 ( rdata_i[10]             ),
       .raddr_o                 ( raddr_o[10]             ),
       .wcoarse_i               ( wcoarse_i[10]           ),
       .rcoarse_o               ( rcoarse_o[10]           ),
       .m0_axi_awvalid          ( m20_axi_awvalid         ),
       .m0_axi_awready          ( m20_axi_awready         ),
       .m0_axi_awaddr           ( m20_axi_awaddr          ),
       .m0_axi_awlen            ( m20_axi_awlen           ),
       .m0_axi_wvalid           ( m20_axi_wvalid          ),
       .m0_axi_wready           ( m20_axi_wready          ),
       .m0_axi_wdata            ( m20_axi_wdata           ),
       .m0_axi_wstrb            ( m20_axi_wstrb           ),
       .m0_axi_wlast            ( m20_axi_wlast           ),
       .m0_axi_bvalid           ( m20_axi_bvalid          ),
       .m0_axi_bready           ( m20_axi_bready          ),
       .m1_axi_awvalid          ( m21_axi_awvalid         ),
       .m1_axi_awready          ( m21_axi_awready         ),
       .m1_axi_awaddr           ( m21_axi_awaddr          ),
       .m1_axi_awlen            ( m21_axi_awlen           ),
       .m1_axi_wvalid           ( m21_axi_wvalid          ),
       .m1_axi_wready           ( m21_axi_wready          ),
       .m1_axi_wdata            ( m21_axi_wdata           ),
       .m1_axi_wstrb            ( m21_axi_wstrb           ),
       .m1_axi_wlast            ( m21_axi_wlast           ),
       .m1_axi_bvalid           ( m21_axi_bvalid          ),
       .m1_axi_bready           ( m21_axi_bready          ),
       .ctrl_addr_offset0       ( axi20_ptr0              ),
       .ctrl_addr_offset1       ( axi21_ptr0              ),
       .dbg_wbeat               (                         ),
       .dbg_wstep               ( dbg_wstep[10]           )
       );

  point_dma_r_channel
    #(
      .ID(22),
      .C_M_AXI_ADDR_WIDTH ( C_M22_AXI_ADDR_WIDTH ),
      .C_M_AXI_DATA_WIDTH ( C_M22_AXI_DATA_WIDTH )
      ) _channel22
      (
       .clk_i,
       .rst_ni,
       .start_i                 ( local_start[22]         ),
       .done_o                  ( local_done[22]          ),
       .hold_o                  ( local_hold[22]          ),
       .release_i               ( local_release[22]       ),
       .we_o                    ( we_o[11]                ),
       .wdata_o                 ( wdata_o[11]             ),
       .waddr_o                 ( waddr_o[11]             ),
       .wcoarse_o               ( wcoarse_o[11]           ),
       .rcoarse_i               ( rcoarse_i[11]           ),
       .m0_axi_arvalid          ( m22_axi_arvalid         ),
       .m0_axi_arready          ( m22_axi_arready         ),
       .m0_axi_araddr           ( m22_axi_araddr          ),
       .m0_axi_arlen            ( m22_axi_arlen           ),
       .m0_axi_rvalid           ( m22_axi_rvalid          ),
       .m0_axi_rready           ( m22_axi_rready          ),
       .m0_axi_rdata            ( m22_axi_rdata           ),
       .m0_axi_rlast            ( m22_axi_rlast           ),
       .m1_axi_arvalid          ( m23_axi_arvalid         ),
       .m1_axi_arready          ( m23_axi_arready         ),
       .m1_axi_araddr           ( m23_axi_araddr          ),
       .m1_axi_arlen            ( m23_axi_arlen           ),
       .m1_axi_rvalid           ( m23_axi_rvalid          ),
       .m1_axi_rready           ( m23_axi_rready          ),
       .m1_axi_rdata            ( m23_axi_rdata           ),
       .m1_axi_rlast            ( m23_axi_rlast           ),
       .ctrl_addr_offset0       ( axi22_ptr0              ),
       .ctrl_addr_offset1       ( axi23_ptr0              ),
       .dbg_rbeat               (                         ),
       .dbg_rstep               ( dbg_rstep[11]           )
       );

  point_dma_w_channel
    #(
      .ID(23),
      .C_M_AXI_ADDR_WIDTH ( C_M23_AXI_ADDR_WIDTH ),
      .C_M_AXI_DATA_WIDTH ( C_M23_AXI_DATA_WIDTH )
      ) _channel23
      (
       .clk_i,
       .rst_ni,
       .start_i                 ( local_start[23]         ),
       .done_o                  ( local_done[23]          ),
       .hold_o                  ( local_hold[23]          ),
       .release_i               ( local_release[23]       ),
       .re_o                    ( re_o[11]                ),
       .rdata_i                 ( rdata_i[11]             ),
       .raddr_o                 ( raddr_o[11]             ),
       .wcoarse_i               ( wcoarse_i[11]           ),
       .rcoarse_o               ( rcoarse_o[11]           ),
       .m0_axi_awvalid          ( m22_axi_awvalid         ),
       .m0_axi_awready          ( m22_axi_awready         ),
       .m0_axi_awaddr           ( m22_axi_awaddr          ),
       .m0_axi_awlen            ( m22_axi_awlen           ),
       .m0_axi_wvalid           ( m22_axi_wvalid          ),
       .m0_axi_wready           ( m22_axi_wready          ),
       .m0_axi_wdata            ( m22_axi_wdata           ),
       .m0_axi_wstrb            ( m22_axi_wstrb           ),
       .m0_axi_wlast            ( m22_axi_wlast           ),
       .m0_axi_bvalid           ( m22_axi_bvalid          ),
       .m0_axi_bready           ( m22_axi_bready          ),
       .m1_axi_awvalid          ( m23_axi_awvalid         ),
       .m1_axi_awready          ( m23_axi_awready         ),
       .m1_axi_awaddr           ( m23_axi_awaddr          ),
       .m1_axi_awlen            ( m23_axi_awlen           ),
       .m1_axi_wvalid           ( m23_axi_wvalid          ),
       .m1_axi_wready           ( m23_axi_wready          ),
       .m1_axi_wdata            ( m23_axi_wdata           ),
       .m1_axi_wstrb            ( m23_axi_wstrb           ),
       .m1_axi_wlast            ( m23_axi_wlast           ),
       .m1_axi_bvalid           ( m23_axi_bvalid          ),
       .m1_axi_bready           ( m23_axi_bready          ),
       .ctrl_addr_offset0       ( axi22_ptr0              ),
       .ctrl_addr_offset1       ( axi23_ptr0              ),
       .dbg_wbeat               (                         ),
       .dbg_wstep               ( dbg_wstep[11]           )
       );

  point_dma_r_channel
    #(
      .ID(24),
      .C_M_AXI_ADDR_WIDTH ( C_M24_AXI_ADDR_WIDTH ),
      .C_M_AXI_DATA_WIDTH ( C_M24_AXI_DATA_WIDTH )
      ) _channel24
      (
       .clk_i,
       .rst_ni,
       .start_i                 ( local_start[24]         ),
       .done_o                  ( local_done[24]          ),
       .hold_o                  ( local_hold[24]          ),
       .release_i               ( local_release[24]       ),
       .we_o                    ( we_o[12]                ),
       .wdata_o                 ( wdata_o[12]             ),
       .waddr_o                 ( waddr_o[12]             ),
       .wcoarse_o               ( wcoarse_o[12]           ),
       .rcoarse_i               ( rcoarse_i[12]           ),
       .m0_axi_arvalid          ( m24_axi_arvalid         ),
       .m0_axi_arready          ( m24_axi_arready         ),
       .m0_axi_araddr           ( m24_axi_araddr          ),
       .m0_axi_arlen            ( m24_axi_arlen           ),
       .m0_axi_rvalid           ( m24_axi_rvalid          ),
       .m0_axi_rready           ( m24_axi_rready          ),
       .m0_axi_rdata            ( m24_axi_rdata           ),
       .m0_axi_rlast            ( m24_axi_rlast           ),
       .m1_axi_arvalid          ( m25_axi_arvalid         ),
       .m1_axi_arready          ( m25_axi_arready         ),
       .m1_axi_araddr           ( m25_axi_araddr          ),
       .m1_axi_arlen            ( m25_axi_arlen           ),
       .m1_axi_rvalid           ( m25_axi_rvalid          ),
       .m1_axi_rready           ( m25_axi_rready          ),
       .m1_axi_rdata            ( m25_axi_rdata           ),
       .m1_axi_rlast            ( m25_axi_rlast           ),
       .ctrl_addr_offset0       ( axi24_ptr0              ),
       .ctrl_addr_offset1       ( axi25_ptr0              ),
       .dbg_rbeat               (                         ),
       .dbg_rstep               ( dbg_rstep[12]           )
       );

  point_dma_w_channel
    #(
      .ID(25),
      .C_M_AXI_ADDR_WIDTH ( C_M25_AXI_ADDR_WIDTH ),
      .C_M_AXI_DATA_WIDTH ( C_M25_AXI_DATA_WIDTH )
      ) _channel25
      (
       .clk_i,
       .rst_ni,
       .start_i                 ( local_start[25]         ),
       .done_o                  ( local_done[25]          ),
       .hold_o                  ( local_hold[25]          ),
       .release_i               ( local_release[25]       ),
       .re_o                    ( re_o[12]                ),
       .rdata_i                 ( rdata_i[12]             ),
       .raddr_o                 ( raddr_o[12]             ),
       .wcoarse_i               ( wcoarse_i[12]           ),
       .rcoarse_o               ( rcoarse_o[12]           ),
       .m0_axi_awvalid          ( m24_axi_awvalid         ),
       .m0_axi_awready          ( m24_axi_awready         ),
       .m0_axi_awaddr           ( m24_axi_awaddr          ),
       .m0_axi_awlen            ( m24_axi_awlen           ),
       .m0_axi_wvalid           ( m24_axi_wvalid          ),
       .m0_axi_wready           ( m24_axi_wready          ),
       .m0_axi_wdata            ( m24_axi_wdata           ),
       .m0_axi_wstrb            ( m24_axi_wstrb           ),
       .m0_axi_wlast            ( m24_axi_wlast           ),
       .m0_axi_bvalid           ( m24_axi_bvalid          ),
       .m0_axi_bready           ( m24_axi_bready          ),
       .m1_axi_awvalid          ( m25_axi_awvalid         ),
       .m1_axi_awready          ( m25_axi_awready         ),
       .m1_axi_awaddr           ( m25_axi_awaddr          ),
       .m1_axi_awlen            ( m25_axi_awlen           ),
       .m1_axi_wvalid           ( m25_axi_wvalid          ),
       .m1_axi_wready           ( m25_axi_wready          ),
       .m1_axi_wdata            ( m25_axi_wdata           ),
       .m1_axi_wstrb            ( m25_axi_wstrb           ),
       .m1_axi_wlast            ( m25_axi_wlast           ),
       .m1_axi_bvalid           ( m25_axi_bvalid          ),
       .m1_axi_bready           ( m25_axi_bready          ),
       .ctrl_addr_offset0       ( axi24_ptr0              ),
       .ctrl_addr_offset1       ( axi25_ptr0              ),
       .dbg_wbeat               (                         ),
       .dbg_wstep               ( dbg_wstep[12]           )
       );

  point_dma_r_channel
    #(
      .ID(26),
      .C_M_AXI_ADDR_WIDTH ( C_M26_AXI_ADDR_WIDTH ),
      .C_M_AXI_DATA_WIDTH ( C_M26_AXI_DATA_WIDTH )
      ) _channel26
      (
       .clk_i,
       .rst_ni,
       .start_i                 ( local_start[26]         ),
       .done_o                  ( local_done[26]          ),
       .hold_o                  ( local_hold[26]          ),
       .release_i               ( local_release[26]       ),
       .we_o                    ( we_o[13]                ),
       .wdata_o                 ( wdata_o[13]             ),
       .waddr_o                 ( waddr_o[13]             ),
       .wcoarse_o               ( wcoarse_o[13]           ),
       .rcoarse_i               ( rcoarse_i[13]           ),
       .m0_axi_arvalid          ( m26_axi_arvalid         ),
       .m0_axi_arready          ( m26_axi_arready         ),
       .m0_axi_araddr           ( m26_axi_araddr          ),
       .m0_axi_arlen            ( m26_axi_arlen           ),
       .m0_axi_rvalid           ( m26_axi_rvalid          ),
       .m0_axi_rready           ( m26_axi_rready          ),
       .m0_axi_rdata            ( m26_axi_rdata           ),
       .m0_axi_rlast            ( m26_axi_rlast           ),
       .m1_axi_arvalid          ( m27_axi_arvalid         ),
       .m1_axi_arready          ( m27_axi_arready         ),
       .m1_axi_araddr           ( m27_axi_araddr          ),
       .m1_axi_arlen            ( m27_axi_arlen           ),
       .m1_axi_rvalid           ( m27_axi_rvalid          ),
       .m1_axi_rready           ( m27_axi_rready          ),
       .m1_axi_rdata            ( m27_axi_rdata           ),
       .m1_axi_rlast            ( m27_axi_rlast           ),
       .ctrl_addr_offset0       ( axi26_ptr0              ),
       .ctrl_addr_offset1       ( axi27_ptr0              ),
       .dbg_rbeat               (                         ),
       .dbg_rstep               ( dbg_rstep[13]           )
       );

  point_dma_w_channel
    #(
      .ID(27),
      .C_M_AXI_ADDR_WIDTH ( C_M27_AXI_ADDR_WIDTH ),
      .C_M_AXI_DATA_WIDTH ( C_M27_AXI_DATA_WIDTH )
      ) _channel27
      (
       .clk_i,
       .rst_ni,
       .start_i                 ( local_start[27]         ),
       .done_o                  ( local_done[27]          ),
       .hold_o                  ( local_hold[27]          ),
       .release_i               ( local_release[27]       ),
       .re_o                    ( re_o[13]                ),
       .rdata_i                 ( rdata_i[13]             ),
       .raddr_o                 ( raddr_o[13]             ),
       .wcoarse_i               ( wcoarse_i[13]           ),
       .rcoarse_o               ( rcoarse_o[13]           ),
       .m0_axi_awvalid          ( m26_axi_awvalid         ),
       .m0_axi_awready          ( m26_axi_awready         ),
       .m0_axi_awaddr           ( m26_axi_awaddr          ),
       .m0_axi_awlen            ( m26_axi_awlen           ),
       .m0_axi_wvalid           ( m26_axi_wvalid          ),
       .m0_axi_wready           ( m26_axi_wready          ),
       .m0_axi_wdata            ( m26_axi_wdata           ),
       .m0_axi_wstrb            ( m26_axi_wstrb           ),
       .m0_axi_wlast            ( m26_axi_wlast           ),
       .m0_axi_bvalid           ( m26_axi_bvalid          ),
       .m0_axi_bready           ( m26_axi_bready          ),
       .m1_axi_awvalid          ( m27_axi_awvalid         ),
       .m1_axi_awready          ( m27_axi_awready         ),
       .m1_axi_awaddr           ( m27_axi_awaddr          ),
       .m1_axi_awlen            ( m27_axi_awlen           ),
       .m1_axi_wvalid           ( m27_axi_wvalid          ),
       .m1_axi_wready           ( m27_axi_wready          ),
       .m1_axi_wdata            ( m27_axi_wdata           ),
       .m1_axi_wstrb            ( m27_axi_wstrb           ),
       .m1_axi_wlast            ( m27_axi_wlast           ),
       .m1_axi_bvalid           ( m27_axi_bvalid          ),
       .m1_axi_bready           ( m27_axi_bready          ),
       .ctrl_addr_offset0       ( axi26_ptr0              ),
       .ctrl_addr_offset1       ( axi27_ptr0              ),
       .dbg_wbeat               (                         ),
       .dbg_wstep               ( dbg_wstep[13]           )
       );

  point_dma_r_channel
    #(
      .ID(28),
      .C_M_AXI_ADDR_WIDTH ( C_M28_AXI_ADDR_WIDTH ),
      .C_M_AXI_DATA_WIDTH ( C_M28_AXI_DATA_WIDTH )
      ) _channel28
      (
       .clk_i,
       .rst_ni,
       .start_i                 ( local_start[28]         ),
       .done_o                  ( local_done[28]          ),
       .hold_o                  ( local_hold[28]          ),
       .release_i               ( local_release[28]       ),
       .we_o                    ( we_o[14]                ),
       .wdata_o                 ( wdata_o[14]             ),
       .waddr_o                 ( waddr_o[14]             ),
       .wcoarse_o               ( wcoarse_o[14]           ),
       .rcoarse_i               ( rcoarse_i[14]           ),
       .m0_axi_arvalid          ( m28_axi_arvalid         ),
       .m0_axi_arready          ( m28_axi_arready         ),
       .m0_axi_araddr           ( m28_axi_araddr          ),
       .m0_axi_arlen            ( m28_axi_arlen           ),
       .m0_axi_rvalid           ( m28_axi_rvalid          ),
       .m0_axi_rready           ( m28_axi_rready          ),
       .m0_axi_rdata            ( m28_axi_rdata           ),
       .m0_axi_rlast            ( m28_axi_rlast           ),
       .m1_axi_arvalid          ( m29_axi_arvalid         ),
       .m1_axi_arready          ( m29_axi_arready         ),
       .m1_axi_araddr           ( m29_axi_araddr          ),
       .m1_axi_arlen            ( m29_axi_arlen           ),
       .m1_axi_rvalid           ( m29_axi_rvalid          ),
       .m1_axi_rready           ( m29_axi_rready          ),
       .m1_axi_rdata            ( m29_axi_rdata           ),
       .m1_axi_rlast            ( m29_axi_rlast           ),
       .ctrl_addr_offset0       ( axi28_ptr0              ),
       .ctrl_addr_offset1       ( axi29_ptr0              ),
       .dbg_rbeat               (                         ),
       .dbg_rstep               ( dbg_rstep[14]           )
       );

  point_dma_w_channel
    #(
      .ID(29),
      .C_M_AXI_ADDR_WIDTH ( C_M29_AXI_ADDR_WIDTH ),
      .C_M_AXI_DATA_WIDTH ( C_M29_AXI_DATA_WIDTH )
      ) _channel29
      (
       .clk_i,
       .rst_ni,
       .start_i                 ( local_start[29]         ),
       .done_o                  ( local_done[29]          ),
       .hold_o                  ( local_hold[29]          ),
       .release_i               ( local_release[29]       ),
       .re_o                    ( re_o[14]                ),
       .rdata_i                 ( rdata_i[14]             ),
       .raddr_o                 ( raddr_o[14]             ),
       .wcoarse_i               ( wcoarse_i[14]           ),
       .rcoarse_o               ( rcoarse_o[14]           ),
       .m0_axi_awvalid          ( m28_axi_awvalid         ),
       .m0_axi_awready          ( m28_axi_awready         ),
       .m0_axi_awaddr           ( m28_axi_awaddr          ),
       .m0_axi_awlen            ( m28_axi_awlen           ),
       .m0_axi_wvalid           ( m28_axi_wvalid          ),
       .m0_axi_wready           ( m28_axi_wready          ),
       .m0_axi_wdata            ( m28_axi_wdata           ),
       .m0_axi_wstrb            ( m28_axi_wstrb           ),
       .m0_axi_wlast            ( m28_axi_wlast           ),
       .m0_axi_bvalid           ( m28_axi_bvalid          ),
       .m0_axi_bready           ( m28_axi_bready          ),
       .m1_axi_awvalid          ( m29_axi_awvalid         ),
       .m1_axi_awready          ( m29_axi_awready         ),
       .m1_axi_awaddr           ( m29_axi_awaddr          ),
       .m1_axi_awlen            ( m29_axi_awlen           ),
       .m1_axi_wvalid           ( m29_axi_wvalid          ),
       .m1_axi_wready           ( m29_axi_wready          ),
       .m1_axi_wdata            ( m29_axi_wdata           ),
       .m1_axi_wstrb            ( m29_axi_wstrb           ),
       .m1_axi_wlast            ( m29_axi_wlast           ),
       .m1_axi_bvalid           ( m29_axi_bvalid          ),
       .m1_axi_bready           ( m29_axi_bready          ),
       .ctrl_addr_offset0       ( axi28_ptr0              ),
       .ctrl_addr_offset1       ( axi29_ptr0              ),
       .dbg_wbeat               (                         ),
       .dbg_wstep               ( dbg_wstep[14]           )
       );

  point_dma_r_channel
    #(
      .ID(30),
      .C_M_AXI_ADDR_WIDTH ( C_M30_AXI_ADDR_WIDTH ),
      .C_M_AXI_DATA_WIDTH ( C_M30_AXI_DATA_WIDTH )
      ) _channel30
      (
       .clk_i,
       .rst_ni,
       .start_i                 ( local_start[30]         ),
       .done_o                  ( local_done[30]          ),
       .hold_o                  ( local_hold[30]          ),
       .release_i               ( local_release[30]       ),
       .we_o                    ( we_o[15]                ),
       .wdata_o                 ( wdata_o[15]             ),
       .waddr_o                 ( waddr_o[15]             ),
       .wcoarse_o               ( wcoarse_o[15]           ),
       .rcoarse_i               ( rcoarse_i[15]           ),
       .m0_axi_arvalid          ( m30_axi_arvalid         ),
       .m0_axi_arready          ( m30_axi_arready         ),
       .m0_axi_araddr           ( m30_axi_araddr          ),
       .m0_axi_arlen            ( m30_axi_arlen           ),
       .m0_axi_rvalid           ( m30_axi_rvalid          ),
       .m0_axi_rready           ( m30_axi_rready          ),
       .m0_axi_rdata            ( m30_axi_rdata           ),
       .m0_axi_rlast            ( m30_axi_rlast           ),
       .m1_axi_arvalid          ( m31_axi_arvalid         ),
       .m1_axi_arready          ( m31_axi_arready         ),
       .m1_axi_araddr           ( m31_axi_araddr          ),
       .m1_axi_arlen            ( m31_axi_arlen           ),
       .m1_axi_rvalid           ( m31_axi_rvalid          ),
       .m1_axi_rready           ( m31_axi_rready          ),
       .m1_axi_rdata            ( m31_axi_rdata           ),
       .m1_axi_rlast            ( m31_axi_rlast           ),
       .ctrl_addr_offset0       ( axi30_ptr0              ),
       .ctrl_addr_offset1       ( axi31_ptr0              ),
       .dbg_rbeat               (                         ),
       .dbg_rstep               ( dbg_rstep[15]           )
       );

  point_dma_w_channel
    #(
      .ID(31),
      .C_M_AXI_ADDR_WIDTH ( C_M31_AXI_ADDR_WIDTH ),
      .C_M_AXI_DATA_WIDTH ( C_M31_AXI_DATA_WIDTH )
      ) _channel31
      (
       .clk_i,
       .rst_ni,
       .start_i                 ( local_start[31]         ),
       .done_o                  ( local_done[31]          ),
       .hold_o                  ( local_hold[31]          ),
       .release_i               ( local_release[31]       ),
       .re_o                    ( re_o[15]                ),
       .rdata_i                 ( rdata_i[15]             ),
       .raddr_o                 ( raddr_o[15]             ),
       .wcoarse_i               ( wcoarse_i[15]           ),
       .rcoarse_o               ( rcoarse_o[15]           ),
       .m0_axi_awvalid          ( m30_axi_awvalid         ),
       .m0_axi_awready          ( m30_axi_awready         ),
       .m0_axi_awaddr           ( m30_axi_awaddr          ),
       .m0_axi_awlen            ( m30_axi_awlen           ),
       .m0_axi_wvalid           ( m30_axi_wvalid          ),
       .m0_axi_wready           ( m30_axi_wready          ),
       .m0_axi_wdata            ( m30_axi_wdata           ),
       .m0_axi_wstrb            ( m30_axi_wstrb           ),
       .m0_axi_wlast            ( m30_axi_wlast           ),
       .m0_axi_bvalid           ( m30_axi_bvalid          ),
       .m0_axi_bready           ( m30_axi_bready          ),
       .m1_axi_awvalid          ( m31_axi_awvalid         ),
       .m1_axi_awready          ( m31_axi_awready         ),
       .m1_axi_awaddr           ( m31_axi_awaddr          ),
       .m1_axi_awlen            ( m31_axi_awlen           ),
       .m1_axi_wvalid           ( m31_axi_wvalid          ),
       .m1_axi_wready           ( m31_axi_wready          ),
       .m1_axi_wdata            ( m31_axi_wdata           ),
       .m1_axi_wstrb            ( m31_axi_wstrb           ),
       .m1_axi_wlast            ( m31_axi_wlast           ),
       .m1_axi_bvalid           ( m31_axi_bvalid          ),
       .m1_axi_bready           ( m31_axi_bready          ),
       .ctrl_addr_offset0       ( axi30_ptr0              ),
       .ctrl_addr_offset1       ( axi31_ptr0              ),
       .dbg_wbeat               (                         ),
       .dbg_wstep               ( dbg_wstep[15]           )
       );

endmodule
