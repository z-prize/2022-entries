// Copyright Supranational LLC
// Licensed under the Apache License, Version 2.0, see LICENSE-APACHE 
// or the MIT license, see LICENSE-MIT, at your option.
// SPDX-License-Identifier: Apache-2.0 OR MIT

(* keep_hierarchy = "yes" *) module ntt_twiddle
  import math_pkg::*;
  #(
    parameter NLEVEL     = 12, // number of butterfly levels (2^12 NTT requires 12 levels)
    parameter NLEVEL0    =  0, // number of mini-cgram levels per stage
    parameter NLANE      =  1, // number of lanes to operate in parallel
    parameter PASS1_ONLY =  0, // 0 for pass 0 or 1 via pass1_i, 1 for pass 1 optimized
    parameter BFLYDSP    = 24  // 24, 16, or 12
    )
  (
   input logic                         rst_ni,
   input logic                         clk_i,

   input logic                         pass1_i,

   output logic [NLANE-1:0][1:0][63:0] w_o,
   input logic [NLANE-1:0]             ready_i
   );


  //
  // In response to reset deassertion or a change in the pass1_i input the twiddle generation
  // will begin priming.  Twiddle factors are generated by ROM lookup and multiplications and
  // ultimately placed in per lane FIFOs at the end of the pipeline.  The depth of the FIFOs
  // needs to be as many cycles as it takes to create and deposit a new twiddle in the FIFO
  // once we see that one has been used.
  //

  localparam CENTRAL_LANE = (NLANE==16) ? 8 : 0;

  localparam PIPE_DEPTH_ROM = 3;
  localparam PIPE_DEPTH_FIFOWR = 1;
  localparam IDEAL_FIFO_DEPTH = PIPE_DEPTH_ROM + PIPE_DEPTH_MULRED + PIPE_DEPTH_FIFOWR;
  localparam FIFO_DEPTH = 1 << $clog2((IDEAL_FIFO_DEPTH < 16) ? 16 : IDEAL_FIFO_DEPTH);
  
  (* dont_touch = "true" *) logic      pass1_untimed_q;
  logic                                restart_a_p0q, restart_b_p0q;
  logic                                restart_p1q, restart_p2q;
  logic [$clog2(FIFO_DEPTH):0]         fifo_count_q;
  logic                                active, advance;

  always_ff @(posedge clk_i) begin
    pass1_untimed_q <= pass1_i;
  end

  ntt_twiddle_restart
    ntt_twiddle_restart
      (
       .clk_i,
       .rst_ni,
       .pass1_i,
       .restart_a_p0q_o(restart_a_p0q),
       .restart_b_p0q_o(restart_b_p0q),
       .restart_p1q_o(restart_p1q),
       .restart_p2q_o(restart_p2q)
       );

  always @(posedge clk_i) begin
    if (restart_b_p0q) begin
      fifo_count_q <= 0;
    end
    else begin
      fifo_count_q
        <= fifo_count_q
           + (active ? 1 : 0)
             - (ready_i[CENTRAL_LANE] ? 1 : 0);
    end
  end


  //
  // For pass==1, the twiddles are the same for all lanes and are provided by the ROM rom_wa.  
  // For pass==0, we can create the per lane twiddles required by combining (mul/reduce) the 
  // rom_wa values with per lane factors which are updated every 2^12 NTT.  The ROM rom_wb 
  // provides the initial value and per 2^12 NTT update values for the factors.

  //
  // Implement rom_wb in "gates".
  //

  localparam [9-1:0][63:0] TWIDDLE_ROM_WB_NLEVEL7
    = 
      {
       64'hbf79143ce60ca966,
       64'h1905d02a5c411f4e,
       64'h9d8f2ad78bfed972,
       64'h0653b4801da1c8cf,
       64'hf2c35199959dfcb6,
       64'h1544ef2335d17997,
       64'he0ee099310bba1e2
       };

  localparam [9-1:0][63:0] TWIDDLE_ROM_WB_NLEVEL9
    = 
      {
       64'h9d8f2ad78bfed972,
       64'h0653b4801da1c8cf,
       64'hf2c35199959dfcb6,
       64'h1544ef2335d17997,
       64'he0ee099310bba1e2,
       64'hf6b2cffe2306baac,
       64'h54df9630bf79450e,
       64'habd0a6e8aa3d8a0e,
       64'h81281a7b05f9beac
       };

  localparam [12-1:0][63:0] TWIDDLE_ROM_WB_NLEVEL12
    = 
      {
       64'h1544ef2335d17997,
       64'he0ee099310bba1e2,
       64'hf6b2cffe2306baac,
       64'h54df9630bf79450e,
       64'habd0a6e8aa3d8a0e,
       64'h81281a7b05f9beac,
       64'hfbd41c6b8caa3302,
       64'h30ba2ecd5e93e76d,
       64'hf502aef532322654,
       64'h4b2a18ade67246b5,
       64'hea9d5a1336fbc98b,
       64'h86cdcc31c307e171
       };

  logic [NLEVEL-1:0][63:0]     rom_wb_small;
  assign rom_wb_small = (NLEVEL== 7) ?  TWIDDLE_ROM_WB_NLEVEL7 :
                        (NLEVEL== 9) ?  TWIDDLE_ROM_WB_NLEVEL9 :
                        (NLEVEL==12) ? TWIDDLE_ROM_WB_NLEVEL12 : 0;

  localparam [63:0] M = 64'hffff_ffff_0000_0001;
  logic [NLANE:0][NLEVEL-1:0][63:0] rom_wb;
  always_comb begin
    for(int i=0;i<NLEVEL;i++) begin
      rom_wb[0][i] = 1;
      for(int j=1;j<NLANE+1;j++) begin
        rom_wb[j][i] = {64'h0,rom_wb[j-1][i]} * {64'h0,rom_wb_small[i]} % M;
      end
    end
  end


  //
  // Pipe stage 0.  Build lookup address for rom_wa and compute rom_wb_level
  //

  logic [NLEVEL-1:0]              i_q, j_q;
  logic [NLEVEL-2:0]              rom_wa_addr_p0;
  logic [$clog2(NLEVEL)-1:0]      rom_wb_level_p0;
  
  always_ff @(posedge clk_i) begin
    if (restart_b_p0q) begin
      i_q <= 0;
      j_q <= 0;
    end
    else begin
      if (advance && active) begin
        if ( (i_q + 2) >= (1 << NLEVEL) ) begin
          i_q <= 0;
          if ( (j_q + NLANE) >= (1 << NLEVEL) ) begin
            j_q <= 0;
          end
          else begin
            j_q <= j_q + NLANE;
          end
        end
        else begin
          i_q <= i_q + 2;
        end
      end
    end
  end

  int                             i_in, z, zz_i, zz_j;
  localparam Nhw = 1<<NLEVEL;
  always_comb begin
    // code here mirrors tb.sv
    i_in = j_q * (1 << NLEVEL) + i_q * NLANE;
    zz_i = i_in / 2 / NLANE % (Nhw/2) / (1 << NLEVEL0);
    zz_j = i_in / 2 / NLANE % (Nhw/2) % (1 << NLEVEL0);
    rom_wa_addr_p0 = zz_j * (1<<(NLEVEL-NLEVEL0-1)) + zz_i;
    for(z=NLEVEL-2;!(rom_wa_addr_p0 & (1 << z)) && z>=0;z--);
    rom_wb_level_p0 = NLEVEL-1-z;
  end


  //
  // Pipe stages 1+2.  Lookup from rom_wa.
  //

  logic [1:0][63:0]               rom_wa_dout_p2;
  logic [$clog2(NLEVEL)-1:0]      rom_wb_level_p1q, rom_wb_level_p2q;
  logic                           valid_p1q, valid_p2q;
  logic                           first_p1q, first_p2q;
  
  always_ff @(posedge clk_i) begin
    valid_p1q <= active && !restart_b_p0q;
    valid_p2q <= valid_p1q;
    rom_wb_level_p1q <= rom_wb_level_p0;
    rom_wb_level_p2q <= rom_wb_level_p1q;
    first_p1q <= (i_q==0) && active && !restart_b_p0q;
    first_p2q <= first_p1q;
  end

  xpm_memory_sprom 
    #(
      .ADDR_WIDTH_A(NLEVEL-1), // DECIMAL
      .AUTO_SLEEP_TIME(0), // DECIMAL
      .CASCADE_HEIGHT(0), // DECIMAL
      .ECC_MODE("no_ecc"), // String
      .MEMORY_INIT_FILE( NLEVEL==7  ? "TWIDDLE_ROM_WA0_NLEVEL7.mem" :
                         NLEVEL==9  ? "TWIDDLE_ROM_WA0_NLEVEL9.mem" : 
                         NLEVEL==12 ? "TWIDDLE_ROM_WA0_NLEVEL12.mem" : "" ),
      .MEMORY_INIT_PARAM(""),
      .MEMORY_OPTIMIZATION("true"), // String
      .MEMORY_PRIMITIVE("auto"), // String
      .MEMORY_SIZE(64<<(NLEVEL-1)), // DECIMAL
      .MESSAGE_CONTROL(0), // DECIMAL
      .READ_DATA_WIDTH_A(64), // DECIMAL
      .READ_LATENCY_A(2), // DECIMAL
      .READ_RESET_VALUE_A("0"), // String
      .RST_MODE_A("SYNC"), // String
      .SIM_ASSERT_CHK(0), // DECIMAL; 0=disable simulation messages, 1=enable simulation messages
      .USE_MEM_INIT(1), // DECIMAL
      .USE_MEM_INIT_MMI(0), // DECIMAL
      .WAKEUP_TIME("disable_sleep") // String
      )
  xpm_memory_sprom0
    (
     .dbiterra(),
     .sbiterra(),
     .douta(rom_wa_dout_p2[0]),
     .addra(rom_wa_addr_p0),
     .clka(clk_i),
     .ena(advance),
     .injectdbiterra(1'b0),
     .injectsbiterra(1'b0),
     .regcea(advance),
     .rsta(1'b0),
     .sleep(1'b0)
     );

  xpm_memory_sprom 
    #(
      .ADDR_WIDTH_A(NLEVEL-1), // DECIMAL
      .AUTO_SLEEP_TIME(0), // DECIMAL
      .CASCADE_HEIGHT(0), // DECIMAL
      .ECC_MODE("no_ecc"), // String
      .MEMORY_INIT_FILE( NLEVEL==7  ? "TWIDDLE_ROM_WA1_NLEVEL7.mem" :
                         NLEVEL==9  ? "TWIDDLE_ROM_WA1_NLEVEL9.mem" : 
                         NLEVEL==12 ? "TWIDDLE_ROM_WA1_NLEVEL12.mem" : "" ),
      .MEMORY_INIT_PARAM(""),
      .MEMORY_OPTIMIZATION("true"), // String
      .MEMORY_PRIMITIVE("auto"), // String
      .MEMORY_SIZE(64<<(NLEVEL-1)), // DECIMAL
      .MESSAGE_CONTROL(0), // DECIMAL
      .READ_DATA_WIDTH_A(64), // DECIMAL
      .READ_LATENCY_A(2), // DECIMAL
      .READ_RESET_VALUE_A("0"), // String
      .RST_MODE_A("SYNC"), // String
      .SIM_ASSERT_CHK(0), // DECIMAL; 0=disable simulation messages, 1=enable simulation messages
      .USE_MEM_INIT(1), // DECIMAL
      .USE_MEM_INIT_MMI(0), // DECIMAL
      .WAKEUP_TIME("disable_sleep") // String
      )
  xpm_memory_sprom1
    (
     .dbiterra(),
     .sbiterra(),
     .douta(rom_wa_dout_p2[1]),
     .addra(rom_wa_addr_p0),
     .clka(clk_i),
     .ena(advance),
     .injectdbiterra(1'b0),
     .injectsbiterra(1'b0),
     .regcea(advance),
     .rsta(1'b0),
     .sleep(1'b0)
     );


  //
  // The below logic is replicated per lane, and will be located near the beginning 
  // of each lane's calculation pipeline.
  //

  if (PASS1_ONLY) begin

    for (genvar gv_i=0; gv_i < NLANE; gv_i++) begin
      assign w_o[gv_i][0] = rom_wa_dout_p2[0];
      assign w_o[gv_i][1] = rom_wa_dout_p2[1];
    end

    assign advance = ready_i[0] || !valid_p2q;
    assign active = 1'b1;

  end

  else begin : pass01


    logic [1:0][63:0] rom_wa_dout_p3q;
  
    always_ff @(posedge clk_i) begin
      rom_wa_dout_p3q <= rom_wa_dout_p2;
    end

    for (genvar gv_i=0; gv_i < NLANE; gv_i++) begin : lane

        ntt_twiddle_lane 
          #(
            .NLEVEL(NLEVEL),
            .BFLYDSP(BFLYDSP), 
            .FIFO_DEPTH(FIFO_DEPTH)
            ) 
        ntt_twiddle_lane
           ( 
             .clk_i,
             .rst_ni,
             .pass1_i,
             .pass1_untimed_i(pass1_untimed_q),
             .first_p2q(first_p2q),
             .valid_p2q(valid_p2q),
             .rom_wb_level_p2q(rom_wb_level_p2q),
             .rom_wb(rom_wb[gv_i]),
             .rom_wb_nlane(rom_wb[NLANE]),
             .rom_wa_dout_p3q(rom_wa_dout_p3q),
             .w_o(w_o[gv_i]),
             .ready_i(ready_i[gv_i])
             );
      
    end

    assign advance = 1'b1;
    assign active = fifo_count_q < FIFO_DEPTH;

  end

endmodule



(* keep_hierarchy = "yes" *) module ntt_twiddle_lane
  import math_pkg::*;
  #(
    parameter NLEVEL = 12,
    parameter BFLYDSP = 24,
    parameter FIFO_DEPTH = 16
    )
  (
   input logic                      clk_i,
   input logic                      rst_ni,
   input logic                      pass1_i,
   input logic                      pass1_untimed_i,
   input logic                      first_p2q,
   input logic                      valid_p2q,
   input logic [$clog2(NLEVEL)-1:0] rom_wb_level_p2q,
   input logic [NLEVEL-1:0][63:0]   rom_wb,
   input logic [NLEVEL-1:0][63:0]   rom_wb_nlane,
   input logic [1:0][63:0]          rom_wa_dout_p3q,
   output logic [1:0][63:0]         w_o,
   input logic                      ready_i
   );
  
  logic                             restart_a_p0q, restart_b_p0q;
  logic                             restart_p1q, restart_p2q;
  
  ntt_twiddle_restart
    ntt_twiddle_restart
      (
       .clk_i,
       .rst_ni,
       .pass1_i,
       .restart_a_p0q_o(restart_a_p0q),
       .restart_b_p0q_o(restart_b_p0q),
       .restart_p1q_o(restart_p1q),
       .restart_p2q_o(restart_p2q)
       );

  //
  // While we are delivering twiddles for the 2^12 NTTs generate the next wb_q 
  // values to use for the next set of NTTs.
  //

  //                   |      |      |      |      |      |      |      |      |
  // restart_a_p0q     |______/-------------\__________________________________________
  // restart_b_p0q     |______/---------------------------\____________________________
  // first_p2q         |xxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx______/------\______________
  // calc_valid_q[0]   |xxxxxxxxxxxxxxxxxxxx\______/--------------------\______________
  // calc_wb_q         |xxxxxxxxxxxxxxxxxxxxxxxxxxx<     rom_wb                ><

  logic [PIPE_DEPTH_MULRED+NLEVEL-1:0] calc_valid_q;
  logic [NLEVEL-1:0][63:0]             calc_wb_q, calc_wb_d;
  logic [63:0]                         calc_w;
  logic [$clog2(NLEVEL)-1:0]           calc_level_q;
  
  always_ff @(posedge clk_i) begin

    if (restart_a_p0q && restart_b_p0q)
      calc_valid_q <= 0;
    else if (!restart_a_p0q && restart_b_p0q)
      calc_valid_q <= 1;
    else if (first_p2q)
      calc_valid_q <= 0;
    else if (!calc_valid_q[0])
      calc_valid_q <= {1'b1,calc_valid_q} >> 1;

    if (restart_b_p0q || first_p2q) begin
      calc_level_q <= 0;
    end
    else if (!calc_valid_q[0]) begin
      calc_level_q <= (calc_level_q==(NLEVEL-1)) ? 0 : (calc_level_q + 1);
    end

  end

  always_comb calc_wb_d = {calc_w, calc_wb_q} >> 64;
  always_ff @(posedge clk_i) begin
    if (!calc_valid_q[0]) begin
      calc_wb_q <= restart_b_p0q ? rom_wb : calc_wb_d;
    end
  end

  mulred #(.BFLYDSP(BFLYDSP)) 
  calc_mulred
    ( .rst_ni(1'b1),
      .clk_i,
      .ce_i(1'b1),
      .a_i(calc_wb_q[0]),
      .b_i(rom_wb_nlane[calc_level_q]),
      .r_o(calc_w)
      );

  //
  // Snapshot the generated wb twiddles when a new 2^12 NTT starts
  //

  logic [NLEVEL-1:0][63:0]          wb_q;
  logic [63:0]                      wb0_q;
  logic                             fifo_rd_ready, fifo_rd_empty, wo_valid_q;
  logic [1:0][63:0]                 w;
  logic [PIPE_DEPTH_MULRED-1:0]     valid_q;     

  always_ff @(posedge clk_i) begin
    if (first_p2q) begin
      wb_q <= calc_wb_q;
    end
    wb0_q <= first_p2q ? 64'h1 : wb_q[rom_wb_level_p2q];
  end
  

  //
  // Perform the multiply and reduction to combine the wa and wb twiddles.
  //

  logic valid_p3q;
  always_ff @(posedge clk_i) begin
    valid_p3q <= valid_p2q;
    valid_q <= restart_p2q ? 0 : ({valid_p3q,valid_q} >> 1);
  end

  mulred #(.BFLYDSP(BFLYDSP)) 
  mulred0
    ( .rst_ni(1'b1),
      .clk_i,
      .ce_i(1'b1),
      .a_i(rom_wa_dout_p3q[0]),
      .b_i(pass1_i ? 64'h1 : wb0_q),
      .r_o(w[0])
      );
  
  mulred #(.BFLYDSP(BFLYDSP)) 
  mulred1
    ( .rst_ni(1'b1),
      .clk_i,
      .ce_i(1'b1),
      .a_i(rom_wa_dout_p3q[1]),
      .b_i(pass1_i ? 64'h1 : wb_q[0]),
      .r_o(w[1])
      );
  
  //
  // Accumulate the generated twiddles in a FIFO and match them up with points when
  // the ready_i signal asserts.
  //

  xpm_fifo_sync 
    #(
      .FIFO_MEMORY_TYPE          ("auto"),                      //string; "auto", "block", "distributed", or "ultra";
      .ECC_MODE                  ("no_ecc"),                    //string; "no_ecc" or "en_ecc";
      .FIFO_WRITE_DEPTH          (FIFO_DEPTH),                  //positive integer
      .WRITE_DATA_WIDTH          (2*64),
      .WR_DATA_COUNT_WIDTH       ($clog2(FIFO_DEPTH)+1),        //positive integer
      .PROG_FULL_THRESH          (10),                          //positive integer, not used
      .FULL_RESET_VALUE          (0),                           //positive integer; 0 or 1
      .READ_MODE                 ("std"),                       //string; "std" or "fwft";
      .FIFO_READ_LATENCY         (1),                           //positive integer;
      .READ_DATA_WIDTH           (2*64),
      .RD_DATA_COUNT_WIDTH       ($clog2(FIFO_DEPTH)+1),
      .PROG_EMPTY_THRESH         (10),                          //positive integer, not used 
      .DOUT_RESET_VALUE          ("0"),                         //string, don't care
      .WAKEUP_TIME               (0)                            //positive integer; 0 or 2;
      ) xpm_fifo_sync
      (
       .sleep         ( 1'b0          ),
       .rst           ( restart_p2q   ),
       .wr_clk        ( clk_i         ),
       .wr_en         ( valid_q[0]    ),
       .din           ( w             ),
       .full          (               ),
       .prog_full     (               ),
       .wr_data_count (               ),
       .overflow      (               ),
       .wr_rst_busy   (               ),
       .almost_full   (               ),
       .wr_ack        (               ),
       .rd_en         ( fifo_rd_ready ),
       .dout          ( w_o           ),
       .empty         ( fifo_rd_empty ),
       .prog_empty    (               ),
       .rd_data_count (               ),
       .underflow     (               ),
       .rd_rst_busy   (               ),
       .almost_empty  (               ),
       .data_valid    (               ),
       .injectsbiterr ( 1'b0          ),
       .injectdbiterr ( 1'b0          ),
       .sbiterr       (               ),
       .dbiterr       (               ) 
       );
  
  assign fifo_rd_ready = !fifo_rd_empty && (!wo_valid_q || ready_i);
  
  always @(posedge clk_i) begin
    if (restart_p2q) begin
      wo_valid_q <= 0;
    end
    else begin
      if (fifo_rd_ready) begin
	wo_valid_q <= 1;
      end
      else if (ready_i) begin
	wo_valid_q <= 0;
      end
    end
  end
  
endmodule


module ntt_twiddle_restart
  #(
    parameter NLEVEL     = 12, // number of butterfly levels (2^12 NTT requires 12 levels)
    parameter NLEVEL0    =  0, // number of mini-cgram levels per stage
    parameter NLANE      =  1, // number of lanes to operate in parallel
    parameter PASS1_ONLY =  0, // 0 for pass 0 or 1 via pass1_i, 1 for pass 1 optimized
    parameter BFLYDSP    = 24  // 24, 16, or 12
    )
  (
   input logic  rst_ni,
   input logic  clk_i,

   input logic  pass1_i,
   output logic restart_a_p0q_o,
   output logic restart_b_p0q_o,
   output logic restart_p1q_o,
   output logic restart_p2q_o
   );

  logic         rst_nq;
  logic [1:0]   pass1_q;
  logic [3:0]   restart_a_p0q, restart_b_p0q;

  always_ff @(posedge clk_i) begin
    rst_nq <= rst_ni;
    pass1_q <= {pass1_q,pass1_i};
  end

  always_ff @(posedge clk_i) begin
    if (!rst_nq || ^pass1_q) begin
      restart_a_p0q <= 4'b0011;
      restart_b_p0q <= 4'b1111;
    end
    else begin
      restart_a_p0q <= restart_a_p0q >> 1;
      restart_b_p0q <= restart_b_p0q >> 1;
    end
  end

  assign restart_a_p0q_o = restart_a_p0q[0];
  assign restart_b_p0q_o = restart_b_p0q[0];

  always_ff @(posedge clk_i) begin
    restart_p1q_o <= restart_b_p0q_o;
    restart_p2q_o <= restart_p1q_o;
  end

endmodule
