// Copyright Supranational LLC
// Licensed under the Apache License, Version 2.0, see LICENSE-APACHE 
// or the MIT license, see LICENSE-MIT, at your option.
// SPDX-License-Identifier: Apache-2.0 OR MIT

// Breaking naming conventions here a bit to speed up
// coding.  Use names that match port names so the
// port wildcarding works.

module nantucket
  #(
    parameter integer C_S_AXI_CONTROL_ADDR_WIDTH = 12 ,
    parameter integer C_S_AXI_CONTROL_DATA_WIDTH = 32 ,
    parameter integer C_M00_AXI_ADDR_WIDTH       = 64 ,
    parameter integer C_M00_AXI_DATA_WIDTH       = 256,
    parameter integer C_M01_AXI_ADDR_WIDTH       = 64 ,
    parameter integer C_M01_AXI_DATA_WIDTH       = 256,
    parameter integer C_M02_AXI_ADDR_WIDTH       = 64 ,
    parameter integer C_M02_AXI_DATA_WIDTH       = 256,
    parameter integer C_M03_AXI_ADDR_WIDTH       = 64 ,
    parameter integer C_M03_AXI_DATA_WIDTH       = 256,
    parameter integer C_M04_AXI_ADDR_WIDTH       = 64 ,
    parameter integer C_M04_AXI_DATA_WIDTH       = 256,
    parameter integer C_M05_AXI_ADDR_WIDTH       = 64 ,
    parameter integer C_M05_AXI_DATA_WIDTH       = 256,
    parameter integer C_M06_AXI_ADDR_WIDTH       = 64 ,
    parameter integer C_M06_AXI_DATA_WIDTH       = 256,
    parameter integer C_M07_AXI_ADDR_WIDTH       = 64 ,
    parameter integer C_M07_AXI_DATA_WIDTH       = 256,
    parameter integer C_M08_AXI_ADDR_WIDTH       = 64 ,
    parameter integer C_M08_AXI_DATA_WIDTH       = 256,
    parameter integer C_M09_AXI_ADDR_WIDTH       = 64 ,
    parameter integer C_M09_AXI_DATA_WIDTH       = 256,
    parameter integer C_M10_AXI_ADDR_WIDTH       = 64 ,
    parameter integer C_M10_AXI_DATA_WIDTH       = 256,
    parameter integer C_M11_AXI_ADDR_WIDTH       = 64 ,
    parameter integer C_M11_AXI_DATA_WIDTH       = 256,
    parameter integer C_M12_AXI_ADDR_WIDTH       = 64 ,
    parameter integer C_M12_AXI_DATA_WIDTH       = 256,
    parameter integer C_M13_AXI_ADDR_WIDTH       = 64 ,
    parameter integer C_M13_AXI_DATA_WIDTH       = 256,
    parameter integer C_M14_AXI_ADDR_WIDTH       = 64 ,
    parameter integer C_M14_AXI_DATA_WIDTH       = 256,
    parameter integer C_M15_AXI_ADDR_WIDTH       = 64 ,
    parameter integer C_M15_AXI_DATA_WIDTH       = 256,
    parameter integer C_M16_AXI_ADDR_WIDTH       = 64 ,
    parameter integer C_M16_AXI_DATA_WIDTH       = 256,
    parameter integer C_M17_AXI_ADDR_WIDTH       = 64 ,
    parameter integer C_M17_AXI_DATA_WIDTH       = 256,
    parameter integer C_M18_AXI_ADDR_WIDTH       = 64 ,
    parameter integer C_M18_AXI_DATA_WIDTH       = 256,
    parameter integer C_M19_AXI_ADDR_WIDTH       = 64 ,
    parameter integer C_M19_AXI_DATA_WIDTH       = 256,
    parameter integer C_M20_AXI_ADDR_WIDTH       = 64 ,
    parameter integer C_M20_AXI_DATA_WIDTH       = 256,
    parameter integer C_M21_AXI_ADDR_WIDTH       = 64 ,
    parameter integer C_M21_AXI_DATA_WIDTH       = 256,
    parameter integer C_M22_AXI_ADDR_WIDTH       = 64 ,
    parameter integer C_M22_AXI_DATA_WIDTH       = 256,
    parameter integer C_M23_AXI_ADDR_WIDTH       = 64 ,
    parameter integer C_M23_AXI_DATA_WIDTH       = 256,
    parameter integer C_M24_AXI_ADDR_WIDTH       = 64 ,
    parameter integer C_M24_AXI_DATA_WIDTH       = 256,
    parameter integer C_M25_AXI_ADDR_WIDTH       = 64 ,
    parameter integer C_M25_AXI_DATA_WIDTH       = 256,
    parameter integer C_M26_AXI_ADDR_WIDTH       = 64 ,
    parameter integer C_M26_AXI_DATA_WIDTH       = 256,
    parameter integer C_M27_AXI_ADDR_WIDTH       = 64 ,
    parameter integer C_M27_AXI_DATA_WIDTH       = 256,
    parameter integer C_M28_AXI_ADDR_WIDTH       = 64 ,
    parameter integer C_M28_AXI_DATA_WIDTH       = 256,
    parameter integer C_M29_AXI_ADDR_WIDTH       = 64 ,
    parameter integer C_M29_AXI_DATA_WIDTH       = 256,
    parameter integer C_M30_AXI_ADDR_WIDTH       = 64 ,
    parameter integer C_M30_AXI_DATA_WIDTH       = 256,
    parameter integer C_M31_AXI_ADDR_WIDTH       = 64 ,
    parameter integer C_M31_AXI_DATA_WIDTH       = 256
    )
  (
   input  wire ap_clk,
   input  wire ap_rst_n,
   input  wire ap_clk_2,
   input  wire ap_rst_n_2,

   // Tool generated ports.
   output wire                              m00_axi_awvalid,
   input  wire                              m00_axi_awready,
   output wire [C_M00_AXI_ADDR_WIDTH-1:0]   m00_axi_awaddr ,
   output wire [8-1:0]                      m00_axi_awlen  ,
   output wire                              m00_axi_wvalid ,
   input  wire                              m00_axi_wready ,
   output wire [C_M00_AXI_DATA_WIDTH-1:0]   m00_axi_wdata  ,
   output wire [C_M00_AXI_DATA_WIDTH/8-1:0] m00_axi_wstrb  ,
   output wire                              m00_axi_wlast  ,
   input  wire                              m00_axi_bvalid ,
   output wire                              m00_axi_bready ,
   output wire                              m00_axi_arvalid,
   input  wire                              m00_axi_arready,
   output wire [C_M00_AXI_ADDR_WIDTH-1:0]   m00_axi_araddr ,
   output wire [8-1:0]                      m00_axi_arlen  ,
   input  wire                              m00_axi_rvalid ,
   output wire                              m00_axi_rready ,
   input  wire [C_M00_AXI_DATA_WIDTH-1:0]   m00_axi_rdata  ,
   input  wire                              m00_axi_rlast  ,

   output wire                              m01_axi_awvalid,
   input  wire                              m01_axi_awready,
   output wire [C_M01_AXI_ADDR_WIDTH-1:0]   m01_axi_awaddr ,
   output wire [8-1:0]                      m01_axi_awlen  ,
   output wire                              m01_axi_wvalid ,
   input  wire                              m01_axi_wready ,
   output wire [C_M01_AXI_DATA_WIDTH-1:0]   m01_axi_wdata  ,
   output wire [C_M01_AXI_DATA_WIDTH/8-1:0] m01_axi_wstrb  ,
   output wire                              m01_axi_wlast  ,
   input  wire                              m01_axi_bvalid ,
   output wire                              m01_axi_bready ,
   output wire                              m01_axi_arvalid,
   input  wire                              m01_axi_arready,
   output wire [C_M01_AXI_ADDR_WIDTH-1:0]   m01_axi_araddr ,
   output wire [8-1:0]                      m01_axi_arlen  ,
   input  wire                              m01_axi_rvalid ,
   output wire                              m01_axi_rready ,
   input  wire [C_M01_AXI_DATA_WIDTH-1:0]   m01_axi_rdata  ,
   input  wire                              m01_axi_rlast  ,

   output wire                              m02_axi_awvalid,
   input  wire                              m02_axi_awready,
   output wire [C_M02_AXI_ADDR_WIDTH-1:0]   m02_axi_awaddr ,
   output wire [8-1:0]                      m02_axi_awlen  ,
   output wire                              m02_axi_wvalid ,
   input  wire                              m02_axi_wready ,
   output wire [C_M02_AXI_DATA_WIDTH-1:0]   m02_axi_wdata  ,
   output wire [C_M02_AXI_DATA_WIDTH/8-1:0] m02_axi_wstrb  ,
   output wire                              m02_axi_wlast  ,
   input  wire                              m02_axi_bvalid ,
   output wire                              m02_axi_bready ,
   output wire                              m02_axi_arvalid,
   input  wire                              m02_axi_arready,
   output wire [C_M02_AXI_ADDR_WIDTH-1:0]   m02_axi_araddr ,
   output wire [8-1:0]                      m02_axi_arlen  ,
   input  wire                              m02_axi_rvalid ,
   output wire                              m02_axi_rready ,
   input  wire [C_M02_AXI_DATA_WIDTH-1:0]   m02_axi_rdata  ,
   input  wire                              m02_axi_rlast  ,

   output wire                              m03_axi_awvalid,
   input  wire                              m03_axi_awready,
   output wire [C_M03_AXI_ADDR_WIDTH-1:0]   m03_axi_awaddr ,
   output wire [8-1:0]                      m03_axi_awlen  ,
   output wire                              m03_axi_wvalid ,
   input  wire                              m03_axi_wready ,
   output wire [C_M03_AXI_DATA_WIDTH-1:0]   m03_axi_wdata  ,
   output wire [C_M03_AXI_DATA_WIDTH/8-1:0] m03_axi_wstrb  ,
   output wire                              m03_axi_wlast  ,
   input  wire                              m03_axi_bvalid ,
   output wire                              m03_axi_bready ,
   output wire                              m03_axi_arvalid,
   input  wire                              m03_axi_arready,
   output wire [C_M03_AXI_ADDR_WIDTH-1:0]   m03_axi_araddr ,
   output wire [8-1:0]                      m03_axi_arlen  ,
   input  wire                              m03_axi_rvalid ,
   output wire                              m03_axi_rready ,
   input  wire [C_M03_AXI_DATA_WIDTH-1:0]   m03_axi_rdata  ,
   input  wire                              m03_axi_rlast  ,

   output wire                              m04_axi_awvalid,
   input  wire                              m04_axi_awready,
   output wire [C_M04_AXI_ADDR_WIDTH-1:0]   m04_axi_awaddr ,
   output wire [8-1:0]                      m04_axi_awlen  ,
   output wire                              m04_axi_wvalid ,
   input  wire                              m04_axi_wready ,
   output wire [C_M04_AXI_DATA_WIDTH-1:0]   m04_axi_wdata  ,
   output wire [C_M04_AXI_DATA_WIDTH/8-1:0] m04_axi_wstrb  ,
   output wire                              m04_axi_wlast  ,
   input  wire                              m04_axi_bvalid ,
   output wire                              m04_axi_bready ,
   output wire                              m04_axi_arvalid,
   input  wire                              m04_axi_arready,
   output wire [C_M04_AXI_ADDR_WIDTH-1:0]   m04_axi_araddr ,
   output wire [8-1:0]                      m04_axi_arlen  ,
   input  wire                              m04_axi_rvalid ,
   output wire                              m04_axi_rready ,
   input  wire [C_M04_AXI_DATA_WIDTH-1:0]   m04_axi_rdata  ,
   input  wire                              m04_axi_rlast  ,

   output wire                              m05_axi_awvalid,
   input  wire                              m05_axi_awready,
   output wire [C_M05_AXI_ADDR_WIDTH-1:0]   m05_axi_awaddr ,
   output wire [8-1:0]                      m05_axi_awlen  ,
   output wire                              m05_axi_wvalid ,
   input  wire                              m05_axi_wready ,
   output wire [C_M05_AXI_DATA_WIDTH-1:0]   m05_axi_wdata  ,
   output wire [C_M05_AXI_DATA_WIDTH/8-1:0] m05_axi_wstrb  ,
   output wire                              m05_axi_wlast  ,
   input  wire                              m05_axi_bvalid ,
   output wire                              m05_axi_bready ,
   output wire                              m05_axi_arvalid,
   input  wire                              m05_axi_arready,
   output wire [C_M05_AXI_ADDR_WIDTH-1:0]   m05_axi_araddr ,
   output wire [8-1:0]                      m05_axi_arlen  ,
   input  wire                              m05_axi_rvalid ,
   output wire                              m05_axi_rready ,
   input  wire [C_M05_AXI_DATA_WIDTH-1:0]   m05_axi_rdata  ,
   input  wire                              m05_axi_rlast  ,

   output wire                              m06_axi_awvalid,
   input  wire                              m06_axi_awready,
   output wire [C_M06_AXI_ADDR_WIDTH-1:0]   m06_axi_awaddr ,
   output wire [8-1:0]                      m06_axi_awlen  ,
   output wire                              m06_axi_wvalid ,
   input  wire                              m06_axi_wready ,
   output wire [C_M06_AXI_DATA_WIDTH-1:0]   m06_axi_wdata  ,
   output wire [C_M06_AXI_DATA_WIDTH/8-1:0] m06_axi_wstrb  ,
   output wire                              m06_axi_wlast  ,
   input  wire                              m06_axi_bvalid ,
   output wire                              m06_axi_bready ,
   output wire                              m06_axi_arvalid,
   input  wire                              m06_axi_arready,
   output wire [C_M06_AXI_ADDR_WIDTH-1:0]   m06_axi_araddr ,
   output wire [8-1:0]                      m06_axi_arlen  ,
   input  wire                              m06_axi_rvalid ,
   output wire                              m06_axi_rready ,
   input  wire [C_M06_AXI_DATA_WIDTH-1:0]   m06_axi_rdata  ,
   input  wire                              m06_axi_rlast  ,

   output wire                              m07_axi_awvalid,
   input  wire                              m07_axi_awready,
   output wire [C_M07_AXI_ADDR_WIDTH-1:0]   m07_axi_awaddr ,
   output wire [8-1:0]                      m07_axi_awlen  ,
   output wire                              m07_axi_wvalid ,
   input  wire                              m07_axi_wready ,
   output wire [C_M07_AXI_DATA_WIDTH-1:0]   m07_axi_wdata  ,
   output wire [C_M07_AXI_DATA_WIDTH/8-1:0] m07_axi_wstrb  ,
   output wire                              m07_axi_wlast  ,
   input  wire                              m07_axi_bvalid ,
   output wire                              m07_axi_bready ,
   output wire                              m07_axi_arvalid,
   input  wire                              m07_axi_arready,
   output wire [C_M07_AXI_ADDR_WIDTH-1:0]   m07_axi_araddr ,
   output wire [8-1:0]                      m07_axi_arlen  ,
   input  wire                              m07_axi_rvalid ,
   output wire                              m07_axi_rready ,
   input  wire [C_M07_AXI_DATA_WIDTH-1:0]   m07_axi_rdata  ,
   input  wire                              m07_axi_rlast  ,

   output wire                              m08_axi_awvalid,
   input  wire                              m08_axi_awready,
   output wire [C_M08_AXI_ADDR_WIDTH-1:0]   m08_axi_awaddr ,
   output wire [8-1:0]                      m08_axi_awlen  ,
   output wire                              m08_axi_wvalid ,
   input  wire                              m08_axi_wready ,
   output wire [C_M08_AXI_DATA_WIDTH-1:0]   m08_axi_wdata  ,
   output wire [C_M08_AXI_DATA_WIDTH/8-1:0] m08_axi_wstrb  ,
   output wire                              m08_axi_wlast  ,
   input  wire                              m08_axi_bvalid ,
   output wire                              m08_axi_bready ,
   output wire                              m08_axi_arvalid,
   input  wire                              m08_axi_arready,
   output wire [C_M08_AXI_ADDR_WIDTH-1:0]   m08_axi_araddr ,
   output wire [8-1:0]                      m08_axi_arlen  ,
   input  wire                              m08_axi_rvalid ,
   output wire                              m08_axi_rready ,
   input  wire [C_M08_AXI_DATA_WIDTH-1:0]   m08_axi_rdata  ,
   input  wire                              m08_axi_rlast  ,

   output wire                              m09_axi_awvalid,
   input  wire                              m09_axi_awready,
   output wire [C_M09_AXI_ADDR_WIDTH-1:0]   m09_axi_awaddr ,
   output wire [8-1:0]                      m09_axi_awlen  ,
   output wire                              m09_axi_wvalid ,
   input  wire                              m09_axi_wready ,
   output wire [C_M09_AXI_DATA_WIDTH-1:0]   m09_axi_wdata  ,
   output wire [C_M09_AXI_DATA_WIDTH/8-1:0] m09_axi_wstrb  ,
   output wire                              m09_axi_wlast  ,
   input  wire                              m09_axi_bvalid ,
   output wire                              m09_axi_bready ,
   output wire                              m09_axi_arvalid,
   input  wire                              m09_axi_arready,
   output wire [C_M09_AXI_ADDR_WIDTH-1:0]   m09_axi_araddr ,
   output wire [8-1:0]                      m09_axi_arlen  ,
   input  wire                              m09_axi_rvalid ,
   output wire                              m09_axi_rready ,
   input  wire [C_M09_AXI_DATA_WIDTH-1:0]   m09_axi_rdata  ,
   input  wire                              m09_axi_rlast  ,

   output wire                              m10_axi_awvalid,
   input  wire                              m10_axi_awready,
   output wire [C_M10_AXI_ADDR_WIDTH-1:0]   m10_axi_awaddr ,
   output wire [8-1:0]                      m10_axi_awlen  ,
   output wire                              m10_axi_wvalid ,
   input  wire                              m10_axi_wready ,
   output wire [C_M10_AXI_DATA_WIDTH-1:0]   m10_axi_wdata  ,
   output wire [C_M10_AXI_DATA_WIDTH/8-1:0] m10_axi_wstrb  ,
   output wire                              m10_axi_wlast  ,
   input  wire                              m10_axi_bvalid ,
   output wire                              m10_axi_bready ,
   output wire                              m10_axi_arvalid,
   input  wire                              m10_axi_arready,
   output wire [C_M10_AXI_ADDR_WIDTH-1:0]   m10_axi_araddr ,
   output wire [8-1:0]                      m10_axi_arlen  ,
   input  wire                              m10_axi_rvalid ,
   output wire                              m10_axi_rready ,
   input  wire [C_M10_AXI_DATA_WIDTH-1:0]   m10_axi_rdata  ,
   input  wire                              m10_axi_rlast  ,

   output wire                              m11_axi_awvalid,
   input  wire                              m11_axi_awready,
   output wire [C_M11_AXI_ADDR_WIDTH-1:0]   m11_axi_awaddr ,
   output wire [8-1:0]                      m11_axi_awlen  ,
   output wire                              m11_axi_wvalid ,
   input  wire                              m11_axi_wready ,
   output wire [C_M11_AXI_DATA_WIDTH-1:0]   m11_axi_wdata  ,
   output wire [C_M11_AXI_DATA_WIDTH/8-1:0] m11_axi_wstrb  ,
   output wire                              m11_axi_wlast  ,
   input  wire                              m11_axi_bvalid ,
   output wire                              m11_axi_bready ,
   output wire                              m11_axi_arvalid,
   input  wire                              m11_axi_arready,
   output wire [C_M11_AXI_ADDR_WIDTH-1:0]   m11_axi_araddr ,
   output wire [8-1:0]                      m11_axi_arlen  ,
   input  wire                              m11_axi_rvalid ,
   output wire                              m11_axi_rready ,
   input  wire [C_M11_AXI_DATA_WIDTH-1:0]   m11_axi_rdata  ,
   input  wire                              m11_axi_rlast  ,

   output wire                              m12_axi_awvalid,
   input  wire                              m12_axi_awready,
   output wire [C_M12_AXI_ADDR_WIDTH-1:0]   m12_axi_awaddr ,
   output wire [8-1:0]                      m12_axi_awlen  ,
   output wire                              m12_axi_wvalid ,
   input  wire                              m12_axi_wready ,
   output wire [C_M12_AXI_DATA_WIDTH-1:0]   m12_axi_wdata  ,
   output wire [C_M12_AXI_DATA_WIDTH/8-1:0] m12_axi_wstrb  ,
   output wire                              m12_axi_wlast  ,
   input  wire                              m12_axi_bvalid ,
   output wire                              m12_axi_bready ,
   output wire                              m12_axi_arvalid,
   input  wire                              m12_axi_arready,
   output wire [C_M12_AXI_ADDR_WIDTH-1:0]   m12_axi_araddr ,
   output wire [8-1:0]                      m12_axi_arlen  ,
   input  wire                              m12_axi_rvalid ,
   output wire                              m12_axi_rready ,
   input  wire [C_M12_AXI_DATA_WIDTH-1:0]   m12_axi_rdata  ,
   input  wire                              m12_axi_rlast  ,

   output wire                              m13_axi_awvalid,
   input  wire                              m13_axi_awready,
   output wire [C_M13_AXI_ADDR_WIDTH-1:0]   m13_axi_awaddr ,
   output wire [8-1:0]                      m13_axi_awlen  ,
   output wire                              m13_axi_wvalid ,
   input  wire                              m13_axi_wready ,
   output wire [C_M13_AXI_DATA_WIDTH-1:0]   m13_axi_wdata  ,
   output wire [C_M13_AXI_DATA_WIDTH/8-1:0] m13_axi_wstrb  ,
   output wire                              m13_axi_wlast  ,
   input  wire                              m13_axi_bvalid ,
   output wire                              m13_axi_bready ,
   output wire                              m13_axi_arvalid,
   input  wire                              m13_axi_arready,
   output wire [C_M13_AXI_ADDR_WIDTH-1:0]   m13_axi_araddr ,
   output wire [8-1:0]                      m13_axi_arlen  ,
   input  wire                              m13_axi_rvalid ,
   output wire                              m13_axi_rready ,
   input  wire [C_M13_AXI_DATA_WIDTH-1:0]   m13_axi_rdata  ,
   input  wire                              m13_axi_rlast  ,

   output wire                              m14_axi_awvalid,
   input  wire                              m14_axi_awready,
   output wire [C_M14_AXI_ADDR_WIDTH-1:0]   m14_axi_awaddr ,
   output wire [8-1:0]                      m14_axi_awlen  ,
   output wire                              m14_axi_wvalid ,
   input  wire                              m14_axi_wready ,
   output wire [C_M14_AXI_DATA_WIDTH-1:0]   m14_axi_wdata  ,
   output wire [C_M14_AXI_DATA_WIDTH/8-1:0] m14_axi_wstrb  ,
   output wire                              m14_axi_wlast  ,
   input  wire                              m14_axi_bvalid ,
   output wire                              m14_axi_bready ,
   output wire                              m14_axi_arvalid,
   input  wire                              m14_axi_arready,
   output wire [C_M14_AXI_ADDR_WIDTH-1:0]   m14_axi_araddr ,
   output wire [8-1:0]                      m14_axi_arlen  ,
   input  wire                              m14_axi_rvalid ,
   output wire                              m14_axi_rready ,
   input  wire [C_M14_AXI_DATA_WIDTH-1:0]   m14_axi_rdata  ,
   input  wire                              m14_axi_rlast  ,

   output wire                              m15_axi_awvalid,
   input  wire                              m15_axi_awready,
   output wire [C_M15_AXI_ADDR_WIDTH-1:0]   m15_axi_awaddr ,
   output wire [8-1:0]                      m15_axi_awlen  ,
   output wire                              m15_axi_wvalid ,
   input  wire                              m15_axi_wready ,
   output wire [C_M15_AXI_DATA_WIDTH-1:0]   m15_axi_wdata  ,
   output wire [C_M15_AXI_DATA_WIDTH/8-1:0] m15_axi_wstrb  ,
   output wire                              m15_axi_wlast  ,
   input  wire                              m15_axi_bvalid ,
   output wire                              m15_axi_bready ,
   output wire                              m15_axi_arvalid,
   input  wire                              m15_axi_arready,
   output wire [C_M15_AXI_ADDR_WIDTH-1:0]   m15_axi_araddr ,
   output wire [8-1:0]                      m15_axi_arlen  ,
   input  wire                              m15_axi_rvalid ,
   output wire                              m15_axi_rready ,
   input  wire [C_M15_AXI_DATA_WIDTH-1:0]   m15_axi_rdata  ,
   input  wire                              m15_axi_rlast  ,

   output wire                              m16_axi_awvalid,
   input  wire                              m16_axi_awready,
   output wire [C_M06_AXI_ADDR_WIDTH-1:0]   m16_axi_awaddr ,
   output wire [8-1:0]                      m16_axi_awlen  ,
   output wire                              m16_axi_wvalid ,
   input  wire                              m16_axi_wready ,
   output wire [C_M06_AXI_DATA_WIDTH-1:0]   m16_axi_wdata  ,
   output wire [C_M06_AXI_DATA_WIDTH/8-1:0] m16_axi_wstrb  ,
   output wire                              m16_axi_wlast  ,
   input  wire                              m16_axi_bvalid ,
   output wire                              m16_axi_bready ,
   output wire                              m16_axi_arvalid,
   input  wire                              m16_axi_arready,
   output wire [C_M06_AXI_ADDR_WIDTH-1:0]   m16_axi_araddr ,
   output wire [8-1:0]                      m16_axi_arlen  ,
   input  wire                              m16_axi_rvalid ,
   output wire                              m16_axi_rready ,
   input  wire [C_M06_AXI_DATA_WIDTH-1:0]   m16_axi_rdata  ,
   input  wire                              m16_axi_rlast  ,

   output wire                              m17_axi_awvalid,
   input  wire                              m17_axi_awready,
   output wire [C_M07_AXI_ADDR_WIDTH-1:0]   m17_axi_awaddr ,
   output wire [8-1:0]                      m17_axi_awlen  ,
   output wire                              m17_axi_wvalid ,
   input  wire                              m17_axi_wready ,
   output wire [C_M07_AXI_DATA_WIDTH-1:0]   m17_axi_wdata  ,
   output wire [C_M07_AXI_DATA_WIDTH/8-1:0] m17_axi_wstrb  ,
   output wire                              m17_axi_wlast  ,
   input  wire                              m17_axi_bvalid ,
   output wire                              m17_axi_bready ,
   output wire                              m17_axi_arvalid,
   input  wire                              m17_axi_arready,
   output wire [C_M07_AXI_ADDR_WIDTH-1:0]   m17_axi_araddr ,
   output wire [8-1:0]                      m17_axi_arlen  ,
   input  wire                              m17_axi_rvalid ,
   output wire                              m17_axi_rready ,
   input  wire [C_M07_AXI_DATA_WIDTH-1:0]   m17_axi_rdata  ,
   input  wire                              m17_axi_rlast  ,

   output wire                              m18_axi_awvalid,
   input  wire                              m18_axi_awready,
   output wire [C_M08_AXI_ADDR_WIDTH-1:0]   m18_axi_awaddr ,
   output wire [8-1:0]                      m18_axi_awlen  ,
   output wire                              m18_axi_wvalid ,
   input  wire                              m18_axi_wready ,
   output wire [C_M08_AXI_DATA_WIDTH-1:0]   m18_axi_wdata  ,
   output wire [C_M08_AXI_DATA_WIDTH/8-1:0] m18_axi_wstrb  ,
   output wire                              m18_axi_wlast  ,
   input  wire                              m18_axi_bvalid ,
   output wire                              m18_axi_bready ,
   output wire                              m18_axi_arvalid,
   input  wire                              m18_axi_arready,
   output wire [C_M08_AXI_ADDR_WIDTH-1:0]   m18_axi_araddr ,
   output wire [8-1:0]                      m18_axi_arlen  ,
   input  wire                              m18_axi_rvalid ,
   output wire                              m18_axi_rready ,
   input  wire [C_M08_AXI_DATA_WIDTH-1:0]   m18_axi_rdata  ,
   input  wire                              m18_axi_rlast  ,

   output wire                              m19_axi_awvalid,
   input  wire                              m19_axi_awready,
   output wire [C_M09_AXI_ADDR_WIDTH-1:0]   m19_axi_awaddr ,
   output wire [8-1:0]                      m19_axi_awlen  ,
   output wire                              m19_axi_wvalid ,
   input  wire                              m19_axi_wready ,
   output wire [C_M09_AXI_DATA_WIDTH-1:0]   m19_axi_wdata  ,
   output wire [C_M09_AXI_DATA_WIDTH/8-1:0] m19_axi_wstrb  ,
   output wire                              m19_axi_wlast  ,
   input  wire                              m19_axi_bvalid ,
   output wire                              m19_axi_bready ,
   output wire                              m19_axi_arvalid,
   input  wire                              m19_axi_arready,
   output wire [C_M09_AXI_ADDR_WIDTH-1:0]   m19_axi_araddr ,
   output wire [8-1:0]                      m19_axi_arlen  ,
   input  wire                              m19_axi_rvalid ,
   output wire                              m19_axi_rready ,
   input  wire [C_M09_AXI_DATA_WIDTH-1:0]   m19_axi_rdata  ,
   input  wire                              m19_axi_rlast  ,

   output wire                              m20_axi_awvalid,
   input  wire                              m20_axi_awready,
   output wire [C_M10_AXI_ADDR_WIDTH-1:0]   m20_axi_awaddr ,
   output wire [8-1:0]                      m20_axi_awlen  ,
   output wire                              m20_axi_wvalid ,
   input  wire                              m20_axi_wready ,
   output wire [C_M10_AXI_DATA_WIDTH-1:0]   m20_axi_wdata  ,
   output wire [C_M10_AXI_DATA_WIDTH/8-1:0] m20_axi_wstrb  ,
   output wire                              m20_axi_wlast  ,
   input  wire                              m20_axi_bvalid ,
   output wire                              m20_axi_bready ,
   output wire                              m20_axi_arvalid,
   input  wire                              m20_axi_arready,
   output wire [C_M10_AXI_ADDR_WIDTH-1:0]   m20_axi_araddr ,
   output wire [8-1:0]                      m20_axi_arlen  ,
   input  wire                              m20_axi_rvalid ,
   output wire                              m20_axi_rready ,
   input  wire [C_M10_AXI_DATA_WIDTH-1:0]   m20_axi_rdata  ,
   input  wire                              m20_axi_rlast  ,

   output wire                              m21_axi_awvalid,
   input  wire                              m21_axi_awready,
   output wire [C_M11_AXI_ADDR_WIDTH-1:0]   m21_axi_awaddr ,
   output wire [8-1:0]                      m21_axi_awlen  ,
   output wire                              m21_axi_wvalid ,
   input  wire                              m21_axi_wready ,
   output wire [C_M11_AXI_DATA_WIDTH-1:0]   m21_axi_wdata  ,
   output wire [C_M11_AXI_DATA_WIDTH/8-1:0] m21_axi_wstrb  ,
   output wire                              m21_axi_wlast  ,
   input  wire                              m21_axi_bvalid ,
   output wire                              m21_axi_bready ,
   output wire                              m21_axi_arvalid,
   input  wire                              m21_axi_arready,
   output wire [C_M11_AXI_ADDR_WIDTH-1:0]   m21_axi_araddr ,
   output wire [8-1:0]                      m21_axi_arlen  ,
   input  wire                              m21_axi_rvalid ,
   output wire                              m21_axi_rready ,
   input  wire [C_M11_AXI_DATA_WIDTH-1:0]   m21_axi_rdata  ,
   input  wire                              m21_axi_rlast  ,

   output wire                              m22_axi_awvalid,
   input  wire                              m22_axi_awready,
   output wire [C_M02_AXI_ADDR_WIDTH-1:0]   m22_axi_awaddr ,
   output wire [8-1:0]                      m22_axi_awlen  ,
   output wire                              m22_axi_wvalid ,
   input  wire                              m22_axi_wready ,
   output wire [C_M02_AXI_DATA_WIDTH-1:0]   m22_axi_wdata  ,
   output wire [C_M02_AXI_DATA_WIDTH/8-1:0] m22_axi_wstrb  ,
   output wire                              m22_axi_wlast  ,
   input  wire                              m22_axi_bvalid ,
   output wire                              m22_axi_bready ,
   output wire                              m22_axi_arvalid,
   input  wire                              m22_axi_arready,
   output wire [C_M02_AXI_ADDR_WIDTH-1:0]   m22_axi_araddr ,
   output wire [8-1:0]                      m22_axi_arlen  ,
   input  wire                              m22_axi_rvalid ,
   output wire                              m22_axi_rready ,
   input  wire [C_M02_AXI_DATA_WIDTH-1:0]   m22_axi_rdata  ,
   input  wire                              m22_axi_rlast  ,

   output wire                              m23_axi_awvalid,
   input  wire                              m23_axi_awready,
   output wire [C_M03_AXI_ADDR_WIDTH-1:0]   m23_axi_awaddr ,
   output wire [8-1:0]                      m23_axi_awlen  ,
   output wire                              m23_axi_wvalid ,
   input  wire                              m23_axi_wready ,
   output wire [C_M03_AXI_DATA_WIDTH-1:0]   m23_axi_wdata  ,
   output wire [C_M03_AXI_DATA_WIDTH/8-1:0] m23_axi_wstrb  ,
   output wire                              m23_axi_wlast  ,
   input  wire                              m23_axi_bvalid ,
   output wire                              m23_axi_bready ,
   output wire                              m23_axi_arvalid,
   input  wire                              m23_axi_arready,
   output wire [C_M03_AXI_ADDR_WIDTH-1:0]   m23_axi_araddr ,
   output wire [8-1:0]                      m23_axi_arlen  ,
   input  wire                              m23_axi_rvalid ,
   output wire                              m23_axi_rready ,
   input  wire [C_M03_AXI_DATA_WIDTH-1:0]   m23_axi_rdata  ,
   input  wire                              m23_axi_rlast  ,

   output wire                              m24_axi_awvalid,
   input  wire                              m24_axi_awready,
   output wire [C_M04_AXI_ADDR_WIDTH-1:0]   m24_axi_awaddr ,
   output wire [8-1:0]                      m24_axi_awlen  ,
   output wire                              m24_axi_wvalid ,
   input  wire                              m24_axi_wready ,
   output wire [C_M04_AXI_DATA_WIDTH-1:0]   m24_axi_wdata  ,
   output wire [C_M04_AXI_DATA_WIDTH/8-1:0] m24_axi_wstrb  ,
   output wire                              m24_axi_wlast  ,
   input  wire                              m24_axi_bvalid ,
   output wire                              m24_axi_bready ,
   output wire                              m24_axi_arvalid,
   input  wire                              m24_axi_arready,
   output wire [C_M04_AXI_ADDR_WIDTH-1:0]   m24_axi_araddr ,
   output wire [8-1:0]                      m24_axi_arlen  ,
   input  wire                              m24_axi_rvalid ,
   output wire                              m24_axi_rready ,
   input  wire [C_M04_AXI_DATA_WIDTH-1:0]   m24_axi_rdata  ,
   input  wire                              m24_axi_rlast  ,

   output wire                              m25_axi_awvalid,
   input  wire                              m25_axi_awready,
   output wire [C_M05_AXI_ADDR_WIDTH-1:0]   m25_axi_awaddr ,
   output wire [8-1:0]                      m25_axi_awlen  ,
   output wire                              m25_axi_wvalid ,
   input  wire                              m25_axi_wready ,
   output wire [C_M05_AXI_DATA_WIDTH-1:0]   m25_axi_wdata  ,
   output wire [C_M05_AXI_DATA_WIDTH/8-1:0] m25_axi_wstrb  ,
   output wire                              m25_axi_wlast  ,
   input  wire                              m25_axi_bvalid ,
   output wire                              m25_axi_bready ,
   output wire                              m25_axi_arvalid,
   input  wire                              m25_axi_arready,
   output wire [C_M05_AXI_ADDR_WIDTH-1:0]   m25_axi_araddr ,
   output wire [8-1:0]                      m25_axi_arlen  ,
   input  wire                              m25_axi_rvalid ,
   output wire                              m25_axi_rready ,
   input  wire [C_M05_AXI_DATA_WIDTH-1:0]   m25_axi_rdata  ,
   input  wire                              m25_axi_rlast  ,

   output wire                              m26_axi_awvalid,
   input  wire                              m26_axi_awready,
   output wire [C_M06_AXI_ADDR_WIDTH-1:0]   m26_axi_awaddr ,
   output wire [8-1:0]                      m26_axi_awlen  ,
   output wire                              m26_axi_wvalid ,
   input  wire                              m26_axi_wready ,
   output wire [C_M06_AXI_DATA_WIDTH-1:0]   m26_axi_wdata  ,
   output wire [C_M06_AXI_DATA_WIDTH/8-1:0] m26_axi_wstrb  ,
   output wire                              m26_axi_wlast  ,
   input  wire                              m26_axi_bvalid ,
   output wire                              m26_axi_bready ,
   output wire                              m26_axi_arvalid,
   input  wire                              m26_axi_arready,
   output wire [C_M06_AXI_ADDR_WIDTH-1:0]   m26_axi_araddr ,
   output wire [8-1:0]                      m26_axi_arlen  ,
   input  wire                              m26_axi_rvalid ,
   output wire                              m26_axi_rready ,
   input  wire [C_M06_AXI_DATA_WIDTH-1:0]   m26_axi_rdata  ,
   input  wire                              m26_axi_rlast  ,

   output wire                              m27_axi_awvalid,
   input  wire                              m27_axi_awready,
   output wire [C_M07_AXI_ADDR_WIDTH-1:0]   m27_axi_awaddr ,
   output wire [8-1:0]                      m27_axi_awlen  ,
   output wire                              m27_axi_wvalid ,
   input  wire                              m27_axi_wready ,
   output wire [C_M07_AXI_DATA_WIDTH-1:0]   m27_axi_wdata  ,
   output wire [C_M07_AXI_DATA_WIDTH/8-1:0] m27_axi_wstrb  ,
   output wire                              m27_axi_wlast  ,
   input  wire                              m27_axi_bvalid ,
   output wire                              m27_axi_bready ,
   output wire                              m27_axi_arvalid,
   input  wire                              m27_axi_arready,
   output wire [C_M07_AXI_ADDR_WIDTH-1:0]   m27_axi_araddr ,
   output wire [8-1:0]                      m27_axi_arlen  ,
   input  wire                              m27_axi_rvalid ,
   output wire                              m27_axi_rready ,
   input  wire [C_M07_AXI_DATA_WIDTH-1:0]   m27_axi_rdata  ,
   input  wire                              m27_axi_rlast  ,

   output wire                              m28_axi_awvalid,
   input  wire                              m28_axi_awready,
   output wire [C_M08_AXI_ADDR_WIDTH-1:0]   m28_axi_awaddr ,
   output wire [8-1:0]                      m28_axi_awlen  ,
   output wire                              m28_axi_wvalid ,
   input  wire                              m28_axi_wready ,
   output wire [C_M08_AXI_DATA_WIDTH-1:0]   m28_axi_wdata  ,
   output wire [C_M08_AXI_DATA_WIDTH/8-1:0] m28_axi_wstrb  ,
   output wire                              m28_axi_wlast  ,
   input  wire                              m28_axi_bvalid ,
   output wire                              m28_axi_bready ,
   output wire                              m28_axi_arvalid,
   input  wire                              m28_axi_arready,
   output wire [C_M08_AXI_ADDR_WIDTH-1:0]   m28_axi_araddr ,
   output wire [8-1:0]                      m28_axi_arlen  ,
   input  wire                              m28_axi_rvalid ,
   output wire                              m28_axi_rready ,
   input  wire [C_M08_AXI_DATA_WIDTH-1:0]   m28_axi_rdata  ,
   input  wire                              m28_axi_rlast  ,

   output wire                              m29_axi_awvalid,
   input  wire                              m29_axi_awready,
   output wire [C_M09_AXI_ADDR_WIDTH-1:0]   m29_axi_awaddr ,
   output wire [8-1:0]                      m29_axi_awlen  ,
   output wire                              m29_axi_wvalid ,
   input  wire                              m29_axi_wready ,
   output wire [C_M09_AXI_DATA_WIDTH-1:0]   m29_axi_wdata  ,
   output wire [C_M09_AXI_DATA_WIDTH/8-1:0] m29_axi_wstrb  ,
   output wire                              m29_axi_wlast  ,
   input  wire                              m29_axi_bvalid ,
   output wire                              m29_axi_bready ,
   output wire                              m29_axi_arvalid,
   input  wire                              m29_axi_arready,
   output wire [C_M09_AXI_ADDR_WIDTH-1:0]   m29_axi_araddr ,
   output wire [8-1:0]                      m29_axi_arlen  ,
   input  wire                              m29_axi_rvalid ,
   output wire                              m29_axi_rready ,
   input  wire [C_M09_AXI_DATA_WIDTH-1:0]   m29_axi_rdata  ,
   input  wire                              m29_axi_rlast  ,

   output wire                              m30_axi_awvalid,
   input  wire                              m30_axi_awready,
   output wire [C_M10_AXI_ADDR_WIDTH-1:0]   m30_axi_awaddr ,
   output wire [8-1:0]                      m30_axi_awlen  ,
   output wire                              m30_axi_wvalid ,
   input  wire                              m30_axi_wready ,
   output wire [C_M10_AXI_DATA_WIDTH-1:0]   m30_axi_wdata  ,
   output wire [C_M10_AXI_DATA_WIDTH/8-1:0] m30_axi_wstrb  ,
   output wire                              m30_axi_wlast  ,
   input  wire                              m30_axi_bvalid ,
   output wire                              m30_axi_bready ,
   output wire                              m30_axi_arvalid,
   input  wire                              m30_axi_arready,
   output wire [C_M10_AXI_ADDR_WIDTH-1:0]   m30_axi_araddr ,
   output wire [8-1:0]                      m30_axi_arlen  ,
   input  wire                              m30_axi_rvalid ,
   output wire                              m30_axi_rready ,
   input  wire [C_M10_AXI_DATA_WIDTH-1:0]   m30_axi_rdata  ,
   input  wire                              m30_axi_rlast  ,

   output wire                              m31_axi_awvalid,
   input  wire                              m31_axi_awready,
   output wire [C_M11_AXI_ADDR_WIDTH-1:0]   m31_axi_awaddr ,
   output wire [8-1:0]                      m31_axi_awlen  ,
   output wire                              m31_axi_wvalid ,
   input  wire                              m31_axi_wready ,
   output wire [C_M11_AXI_DATA_WIDTH-1:0]   m31_axi_wdata  ,
   output wire [C_M11_AXI_DATA_WIDTH/8-1:0] m31_axi_wstrb  ,
   output wire                              m31_axi_wlast  ,
   input  wire                              m31_axi_bvalid ,
   output wire                              m31_axi_bready ,
   output wire                              m31_axi_arvalid,
   input  wire                              m31_axi_arready,
   output wire [C_M11_AXI_ADDR_WIDTH-1:0]   m31_axi_araddr ,
   output wire [8-1:0]                      m31_axi_arlen  ,
   input  wire                              m31_axi_rvalid ,
   output wire                              m31_axi_rready ,
   input  wire [C_M11_AXI_DATA_WIDTH-1:0]   m31_axi_rdata  ,
   input  wire                              m31_axi_rlast  ,

   input  wire                                    s_axi_control_awvalid,
   output wire                                    s_axi_control_awready,
   input  wire [C_S_AXI_CONTROL_ADDR_WIDTH-1:0]   s_axi_control_awaddr ,
   input  wire                                    s_axi_control_wvalid ,
   output wire                                    s_axi_control_wready ,
   input  wire [C_S_AXI_CONTROL_DATA_WIDTH-1:0]   s_axi_control_wdata  ,
   input  wire [C_S_AXI_CONTROL_DATA_WIDTH/8-1:0] s_axi_control_wstrb  ,
   input  wire                                    s_axi_control_arvalid,
   output wire                                    s_axi_control_arready,
   input  wire [C_S_AXI_CONTROL_ADDR_WIDTH-1:0]   s_axi_control_araddr ,
   output wire                                    s_axi_control_rvalid ,
   input  wire                                    s_axi_control_rready ,
   output wire [C_S_AXI_CONTROL_DATA_WIDTH-1:0]   s_axi_control_rdata  ,
   output wire [2-1:0]                            s_axi_control_rresp  ,
   output wire                                    s_axi_control_bvalid ,
   input  wire                                    s_axi_control_bready ,
   output wire [2-1:0]                            s_axi_control_bresp  ,

   output wire                                    interrupt            
   );

  nantucket_sv
    #(
      .C_S_AXI_CONTROL_ADDR_WIDTH ( C_S_AXI_CONTROL_ADDR_WIDTH ),
      .C_S_AXI_CONTROL_DATA_WIDTH ( C_S_AXI_CONTROL_DATA_WIDTH ),
      .C_M00_AXI_ADDR_WIDTH ( C_M00_AXI_ADDR_WIDTH ),
      .C_M00_AXI_DATA_WIDTH ( C_M00_AXI_DATA_WIDTH ),
      .C_M01_AXI_ADDR_WIDTH ( C_M01_AXI_ADDR_WIDTH ),
      .C_M01_AXI_DATA_WIDTH ( C_M01_AXI_DATA_WIDTH ),
      .C_M02_AXI_ADDR_WIDTH ( C_M02_AXI_ADDR_WIDTH ),
      .C_M02_AXI_DATA_WIDTH ( C_M02_AXI_DATA_WIDTH ),
      .C_M03_AXI_ADDR_WIDTH ( C_M03_AXI_ADDR_WIDTH ),
      .C_M03_AXI_DATA_WIDTH ( C_M03_AXI_DATA_WIDTH ),
      .C_M04_AXI_ADDR_WIDTH ( C_M04_AXI_ADDR_WIDTH ),
      .C_M04_AXI_DATA_WIDTH ( C_M04_AXI_DATA_WIDTH ),
      .C_M05_AXI_ADDR_WIDTH ( C_M05_AXI_ADDR_WIDTH ),
      .C_M05_AXI_DATA_WIDTH ( C_M05_AXI_DATA_WIDTH ),
      .C_M06_AXI_ADDR_WIDTH ( C_M06_AXI_ADDR_WIDTH ),
      .C_M06_AXI_DATA_WIDTH ( C_M06_AXI_DATA_WIDTH ),
      .C_M07_AXI_ADDR_WIDTH ( C_M07_AXI_ADDR_WIDTH ),
      .C_M07_AXI_DATA_WIDTH ( C_M07_AXI_DATA_WIDTH ),
      .C_M08_AXI_ADDR_WIDTH ( C_M08_AXI_ADDR_WIDTH ),
      .C_M08_AXI_DATA_WIDTH ( C_M08_AXI_DATA_WIDTH ),
      .C_M09_AXI_ADDR_WIDTH ( C_M09_AXI_ADDR_WIDTH ),
      .C_M09_AXI_DATA_WIDTH ( C_M09_AXI_DATA_WIDTH ),
      .C_M10_AXI_ADDR_WIDTH ( C_M10_AXI_ADDR_WIDTH ),
      .C_M10_AXI_DATA_WIDTH ( C_M10_AXI_DATA_WIDTH ),
      .C_M11_AXI_ADDR_WIDTH ( C_M11_AXI_ADDR_WIDTH ),
      .C_M11_AXI_DATA_WIDTH ( C_M11_AXI_DATA_WIDTH ),
      .C_M12_AXI_ADDR_WIDTH ( C_M12_AXI_ADDR_WIDTH ),
      .C_M12_AXI_DATA_WIDTH ( C_M12_AXI_DATA_WIDTH ),
      .C_M13_AXI_ADDR_WIDTH ( C_M13_AXI_ADDR_WIDTH ),
      .C_M13_AXI_DATA_WIDTH ( C_M13_AXI_DATA_WIDTH ),
      .C_M14_AXI_ADDR_WIDTH ( C_M14_AXI_ADDR_WIDTH ),
      .C_M14_AXI_DATA_WIDTH ( C_M14_AXI_DATA_WIDTH ),
      .C_M15_AXI_ADDR_WIDTH ( C_M15_AXI_ADDR_WIDTH ),
      .C_M15_AXI_DATA_WIDTH ( C_M15_AXI_DATA_WIDTH ),
      .C_M16_AXI_ADDR_WIDTH ( C_M16_AXI_ADDR_WIDTH ),
      .C_M16_AXI_DATA_WIDTH ( C_M16_AXI_DATA_WIDTH ),
      .C_M17_AXI_ADDR_WIDTH ( C_M17_AXI_ADDR_WIDTH ),
      .C_M17_AXI_DATA_WIDTH ( C_M17_AXI_DATA_WIDTH ),
      .C_M18_AXI_ADDR_WIDTH ( C_M18_AXI_ADDR_WIDTH ),
      .C_M18_AXI_DATA_WIDTH ( C_M18_AXI_DATA_WIDTH ),
      .C_M19_AXI_ADDR_WIDTH ( C_M19_AXI_ADDR_WIDTH ),
      .C_M19_AXI_DATA_WIDTH ( C_M19_AXI_DATA_WIDTH ),
      .C_M20_AXI_ADDR_WIDTH ( C_M20_AXI_ADDR_WIDTH ),
      .C_M20_AXI_DATA_WIDTH ( C_M20_AXI_DATA_WIDTH ),
      .C_M21_AXI_ADDR_WIDTH ( C_M21_AXI_ADDR_WIDTH ),
      .C_M21_AXI_DATA_WIDTH ( C_M21_AXI_DATA_WIDTH ),
      .C_M22_AXI_ADDR_WIDTH ( C_M22_AXI_ADDR_WIDTH ),
      .C_M22_AXI_DATA_WIDTH ( C_M22_AXI_DATA_WIDTH ),
      .C_M23_AXI_ADDR_WIDTH ( C_M23_AXI_ADDR_WIDTH ),
      .C_M23_AXI_DATA_WIDTH ( C_M23_AXI_DATA_WIDTH ),
      .C_M24_AXI_ADDR_WIDTH ( C_M24_AXI_ADDR_WIDTH ),
      .C_M24_AXI_DATA_WIDTH ( C_M24_AXI_DATA_WIDTH ),
      .C_M25_AXI_ADDR_WIDTH ( C_M25_AXI_ADDR_WIDTH ),
      .C_M25_AXI_DATA_WIDTH ( C_M25_AXI_DATA_WIDTH ),
      .C_M26_AXI_ADDR_WIDTH ( C_M26_AXI_ADDR_WIDTH ),
      .C_M26_AXI_DATA_WIDTH ( C_M26_AXI_DATA_WIDTH ),
      .C_M27_AXI_ADDR_WIDTH ( C_M27_AXI_ADDR_WIDTH ),
      .C_M27_AXI_DATA_WIDTH ( C_M27_AXI_DATA_WIDTH ),
      .C_M28_AXI_ADDR_WIDTH ( C_M28_AXI_ADDR_WIDTH ),
      .C_M28_AXI_DATA_WIDTH ( C_M28_AXI_DATA_WIDTH ),
      .C_M29_AXI_ADDR_WIDTH ( C_M29_AXI_ADDR_WIDTH ),
      .C_M29_AXI_DATA_WIDTH ( C_M29_AXI_DATA_WIDTH ),
      .C_M30_AXI_ADDR_WIDTH ( C_M30_AXI_ADDR_WIDTH ),
      .C_M30_AXI_DATA_WIDTH ( C_M30_AXI_DATA_WIDTH ),
      .C_M31_AXI_ADDR_WIDTH ( C_M31_AXI_ADDR_WIDTH ),
      .C_M31_AXI_DATA_WIDTH ( C_M31_AXI_DATA_WIDTH )
      ) _nantucket_sv
      (
       .dma_clk_i(ap_clk),
       .dma_rst_ni(ap_rst_n),
       .ntt_clk_i(ap_clk_2),

       .m00_axi_awvalid(m00_axi_awvalid),
       .m00_axi_awready(m00_axi_awready),
       .m00_axi_awaddr(m00_axi_awaddr),
       .m00_axi_awlen(m00_axi_awlen),
       .m00_axi_wvalid(m00_axi_wvalid),
       .m00_axi_wready(m00_axi_wready),
       .m00_axi_wdata(m00_axi_wdata),
       .m00_axi_wstrb(m00_axi_wstrb),
       .m00_axi_wlast(m00_axi_wlast),
       .m00_axi_bvalid(m00_axi_bvalid),
       .m00_axi_bready(m00_axi_bready),
       .m00_axi_arvalid(m00_axi_arvalid),
       .m00_axi_arready(m00_axi_arready),
       .m00_axi_araddr(m00_axi_araddr),
       .m00_axi_arlen(m00_axi_arlen),
       .m00_axi_rvalid(m00_axi_rvalid),
       .m00_axi_rready(m00_axi_rready),
       .m00_axi_rdata(m00_axi_rdata),
       .m00_axi_rlast(m00_axi_rlast),

       .m01_axi_awvalid(m01_axi_awvalid),
       .m01_axi_awready(m01_axi_awready),
       .m01_axi_awaddr(m01_axi_awaddr),
       .m01_axi_awlen(m01_axi_awlen),
       .m01_axi_wvalid(m01_axi_wvalid),
       .m01_axi_wready(m01_axi_wready),
       .m01_axi_wdata(m01_axi_wdata),
       .m01_axi_wstrb(m01_axi_wstrb),
       .m01_axi_wlast(m01_axi_wlast),
       .m01_axi_bvalid(m01_axi_bvalid),
       .m01_axi_bready(m01_axi_bready),
       .m01_axi_arvalid(m01_axi_arvalid),
       .m01_axi_arready(m01_axi_arready),
       .m01_axi_araddr(m01_axi_araddr),
       .m01_axi_arlen(m01_axi_arlen),
       .m01_axi_rvalid(m01_axi_rvalid),
       .m01_axi_rready(m01_axi_rready),
       .m01_axi_rdata(m01_axi_rdata),
       .m01_axi_rlast(m01_axi_rlast),

       .m02_axi_awvalid(m02_axi_awvalid),
       .m02_axi_awready(m02_axi_awready),
       .m02_axi_awaddr(m02_axi_awaddr),
       .m02_axi_awlen(m02_axi_awlen),
       .m02_axi_wvalid(m02_axi_wvalid),
       .m02_axi_wready(m02_axi_wready),
       .m02_axi_wdata(m02_axi_wdata),
       .m02_axi_wstrb(m02_axi_wstrb),
       .m02_axi_wlast(m02_axi_wlast),
       .m02_axi_bvalid(m02_axi_bvalid),
       .m02_axi_bready(m02_axi_bready),
       .m02_axi_arvalid(m02_axi_arvalid),
       .m02_axi_arready(m02_axi_arready),
       .m02_axi_araddr(m02_axi_araddr),
       .m02_axi_arlen(m02_axi_arlen),
       .m02_axi_rvalid(m02_axi_rvalid),
       .m02_axi_rready(m02_axi_rready),
       .m02_axi_rdata(m02_axi_rdata),
       .m02_axi_rlast(m02_axi_rlast),

       .m03_axi_awvalid(m03_axi_awvalid),
       .m03_axi_awready(m03_axi_awready),
       .m03_axi_awaddr(m03_axi_awaddr),
       .m03_axi_awlen(m03_axi_awlen),
       .m03_axi_wvalid(m03_axi_wvalid),
       .m03_axi_wready(m03_axi_wready),
       .m03_axi_wdata(m03_axi_wdata),
       .m03_axi_wstrb(m03_axi_wstrb),
       .m03_axi_wlast(m03_axi_wlast),
       .m03_axi_bvalid(m03_axi_bvalid),
       .m03_axi_bready(m03_axi_bready),
       .m03_axi_arvalid(m03_axi_arvalid),
       .m03_axi_arready(m03_axi_arready),
       .m03_axi_araddr(m03_axi_araddr),
       .m03_axi_arlen(m03_axi_arlen),
       .m03_axi_rvalid(m03_axi_rvalid),
       .m03_axi_rready(m03_axi_rready),
       .m03_axi_rdata(m03_axi_rdata),
       .m03_axi_rlast(m03_axi_rlast),

       .m04_axi_awvalid(m04_axi_awvalid),
       .m04_axi_awready(m04_axi_awready),
       .m04_axi_awaddr(m04_axi_awaddr),
       .m04_axi_awlen(m04_axi_awlen),
       .m04_axi_wvalid(m04_axi_wvalid),
       .m04_axi_wready(m04_axi_wready),
       .m04_axi_wdata(m04_axi_wdata),
       .m04_axi_wstrb(m04_axi_wstrb),
       .m04_axi_wlast(m04_axi_wlast),
       .m04_axi_bvalid(m04_axi_bvalid),
       .m04_axi_bready(m04_axi_bready),
       .m04_axi_arvalid(m04_axi_arvalid),
       .m04_axi_arready(m04_axi_arready),
       .m04_axi_araddr(m04_axi_araddr),
       .m04_axi_arlen(m04_axi_arlen),
       .m04_axi_rvalid(m04_axi_rvalid),
       .m04_axi_rready(m04_axi_rready),
       .m04_axi_rdata(m04_axi_rdata),
       .m04_axi_rlast(m04_axi_rlast),

       .m05_axi_awvalid(m05_axi_awvalid),
       .m05_axi_awready(m05_axi_awready),
       .m05_axi_awaddr(m05_axi_awaddr),
       .m05_axi_awlen(m05_axi_awlen),
       .m05_axi_wvalid(m05_axi_wvalid),
       .m05_axi_wready(m05_axi_wready),
       .m05_axi_wdata(m05_axi_wdata),
       .m05_axi_wstrb(m05_axi_wstrb),
       .m05_axi_wlast(m05_axi_wlast),
       .m05_axi_bvalid(m05_axi_bvalid),
       .m05_axi_bready(m05_axi_bready),
       .m05_axi_arvalid(m05_axi_arvalid),
       .m05_axi_arready(m05_axi_arready),
       .m05_axi_araddr(m05_axi_araddr),
       .m05_axi_arlen(m05_axi_arlen),
       .m05_axi_rvalid(m05_axi_rvalid),
       .m05_axi_rready(m05_axi_rready),
       .m05_axi_rdata(m05_axi_rdata),
       .m05_axi_rlast(m05_axi_rlast),

       .m06_axi_awvalid(m06_axi_awvalid),
       .m06_axi_awready(m06_axi_awready),
       .m06_axi_awaddr(m06_axi_awaddr),
       .m06_axi_awlen(m06_axi_awlen),
       .m06_axi_wvalid(m06_axi_wvalid),
       .m06_axi_wready(m06_axi_wready),
       .m06_axi_wdata(m06_axi_wdata),
       .m06_axi_wstrb(m06_axi_wstrb),
       .m06_axi_wlast(m06_axi_wlast),
       .m06_axi_bvalid(m06_axi_bvalid),
       .m06_axi_bready(m06_axi_bready),
       .m06_axi_arvalid(m06_axi_arvalid),
       .m06_axi_arready(m06_axi_arready),
       .m06_axi_araddr(m06_axi_araddr),
       .m06_axi_arlen(m06_axi_arlen),
       .m06_axi_rvalid(m06_axi_rvalid),
       .m06_axi_rready(m06_axi_rready),
       .m06_axi_rdata(m06_axi_rdata),
       .m06_axi_rlast(m06_axi_rlast),

       .m07_axi_awvalid(m07_axi_awvalid),
       .m07_axi_awready(m07_axi_awready),
       .m07_axi_awaddr(m07_axi_awaddr),
       .m07_axi_awlen(m07_axi_awlen),
       .m07_axi_wvalid(m07_axi_wvalid),
       .m07_axi_wready(m07_axi_wready),
       .m07_axi_wdata(m07_axi_wdata),
       .m07_axi_wstrb(m07_axi_wstrb),
       .m07_axi_wlast(m07_axi_wlast),
       .m07_axi_bvalid(m07_axi_bvalid),
       .m07_axi_bready(m07_axi_bready),
       .m07_axi_arvalid(m07_axi_arvalid),
       .m07_axi_arready(m07_axi_arready),
       .m07_axi_araddr(m07_axi_araddr),
       .m07_axi_arlen(m07_axi_arlen),
       .m07_axi_rvalid(m07_axi_rvalid),
       .m07_axi_rready(m07_axi_rready),
       .m07_axi_rdata(m07_axi_rdata),
       .m07_axi_rlast(m07_axi_rlast),

       .m08_axi_awvalid(m08_axi_awvalid),
       .m08_axi_awready(m08_axi_awready),
       .m08_axi_awaddr(m08_axi_awaddr),
       .m08_axi_awlen(m08_axi_awlen),
       .m08_axi_wvalid(m08_axi_wvalid),
       .m08_axi_wready(m08_axi_wready),
       .m08_axi_wdata(m08_axi_wdata),
       .m08_axi_wstrb(m08_axi_wstrb),
       .m08_axi_wlast(m08_axi_wlast),
       .m08_axi_bvalid(m08_axi_bvalid),
       .m08_axi_bready(m08_axi_bready),
       .m08_axi_arvalid(m08_axi_arvalid),
       .m08_axi_arready(m08_axi_arready),
       .m08_axi_araddr(m08_axi_araddr),
       .m08_axi_arlen(m08_axi_arlen),
       .m08_axi_rvalid(m08_axi_rvalid),
       .m08_axi_rready(m08_axi_rready),
       .m08_axi_rdata(m08_axi_rdata),
       .m08_axi_rlast(m08_axi_rlast),

       .m09_axi_awvalid(m09_axi_awvalid),
       .m09_axi_awready(m09_axi_awready),
       .m09_axi_awaddr(m09_axi_awaddr),
       .m09_axi_awlen(m09_axi_awlen),
       .m09_axi_wvalid(m09_axi_wvalid),
       .m09_axi_wready(m09_axi_wready),
       .m09_axi_wdata(m09_axi_wdata),
       .m09_axi_wstrb(m09_axi_wstrb),
       .m09_axi_wlast(m09_axi_wlast),
       .m09_axi_bvalid(m09_axi_bvalid),
       .m09_axi_bready(m09_axi_bready),
       .m09_axi_arvalid(m09_axi_arvalid),
       .m09_axi_arready(m09_axi_arready),
       .m09_axi_araddr(m09_axi_araddr),
       .m09_axi_arlen(m09_axi_arlen),
       .m09_axi_rvalid(m09_axi_rvalid),
       .m09_axi_rready(m09_axi_rready),
       .m09_axi_rdata(m09_axi_rdata),
       .m09_axi_rlast(m09_axi_rlast),

       .m10_axi_awvalid(m10_axi_awvalid),
       .m10_axi_awready(m10_axi_awready),
       .m10_axi_awaddr(m10_axi_awaddr),
       .m10_axi_awlen(m10_axi_awlen),
       .m10_axi_wvalid(m10_axi_wvalid),
       .m10_axi_wready(m10_axi_wready),
       .m10_axi_wdata(m10_axi_wdata),
       .m10_axi_wstrb(m10_axi_wstrb),
       .m10_axi_wlast(m10_axi_wlast),
       .m10_axi_bvalid(m10_axi_bvalid),
       .m10_axi_bready(m10_axi_bready),
       .m10_axi_arvalid(m10_axi_arvalid),
       .m10_axi_arready(m10_axi_arready),
       .m10_axi_araddr(m10_axi_araddr),
       .m10_axi_arlen(m10_axi_arlen),
       .m10_axi_rvalid(m10_axi_rvalid),
       .m10_axi_rready(m10_axi_rready),
       .m10_axi_rdata(m10_axi_rdata),
       .m10_axi_rlast(m10_axi_rlast),

       .m11_axi_awvalid(m11_axi_awvalid),
       .m11_axi_awready(m11_axi_awready),
       .m11_axi_awaddr(m11_axi_awaddr),
       .m11_axi_awlen(m11_axi_awlen),
       .m11_axi_wvalid(m11_axi_wvalid),
       .m11_axi_wready(m11_axi_wready),
       .m11_axi_wdata(m11_axi_wdata),
       .m11_axi_wstrb(m11_axi_wstrb),
       .m11_axi_wlast(m11_axi_wlast),
       .m11_axi_bvalid(m11_axi_bvalid),
       .m11_axi_bready(m11_axi_bready),
       .m11_axi_arvalid(m11_axi_arvalid),
       .m11_axi_arready(m11_axi_arready),
       .m11_axi_araddr(m11_axi_araddr),
       .m11_axi_arlen(m11_axi_arlen),
       .m11_axi_rvalid(m11_axi_rvalid),
       .m11_axi_rready(m11_axi_rready),
       .m11_axi_rdata(m11_axi_rdata),
       .m11_axi_rlast(m11_axi_rlast),

       .m12_axi_awvalid(m12_axi_awvalid),
       .m12_axi_awready(m12_axi_awready),
       .m12_axi_awaddr(m12_axi_awaddr),
       .m12_axi_awlen(m12_axi_awlen),
       .m12_axi_wvalid(m12_axi_wvalid),
       .m12_axi_wready(m12_axi_wready),
       .m12_axi_wdata(m12_axi_wdata),
       .m12_axi_wstrb(m12_axi_wstrb),
       .m12_axi_wlast(m12_axi_wlast),
       .m12_axi_bvalid(m12_axi_bvalid),
       .m12_axi_bready(m12_axi_bready),
       .m12_axi_arvalid(m12_axi_arvalid),
       .m12_axi_arready(m12_axi_arready),
       .m12_axi_araddr(m12_axi_araddr),
       .m12_axi_arlen(m12_axi_arlen),
       .m12_axi_rvalid(m12_axi_rvalid),
       .m12_axi_rready(m12_axi_rready),
       .m12_axi_rdata(m12_axi_rdata),
       .m12_axi_rlast(m12_axi_rlast),

       .m13_axi_awvalid(m13_axi_awvalid),
       .m13_axi_awready(m13_axi_awready),
       .m13_axi_awaddr(m13_axi_awaddr),
       .m13_axi_awlen(m13_axi_awlen),
       .m13_axi_wvalid(m13_axi_wvalid),
       .m13_axi_wready(m13_axi_wready),
       .m13_axi_wdata(m13_axi_wdata),
       .m13_axi_wstrb(m13_axi_wstrb),
       .m13_axi_wlast(m13_axi_wlast),
       .m13_axi_bvalid(m13_axi_bvalid),
       .m13_axi_bready(m13_axi_bready),
       .m13_axi_arvalid(m13_axi_arvalid),
       .m13_axi_arready(m13_axi_arready),
       .m13_axi_araddr(m13_axi_araddr),
       .m13_axi_arlen(m13_axi_arlen),
       .m13_axi_rvalid(m13_axi_rvalid),
       .m13_axi_rready(m13_axi_rready),
       .m13_axi_rdata(m13_axi_rdata),
       .m13_axi_rlast(m13_axi_rlast),

       .m14_axi_awvalid(m14_axi_awvalid),
       .m14_axi_awready(m14_axi_awready),
       .m14_axi_awaddr(m14_axi_awaddr),
       .m14_axi_awlen(m14_axi_awlen),
       .m14_axi_wvalid(m14_axi_wvalid),
       .m14_axi_wready(m14_axi_wready),
       .m14_axi_wdata(m14_axi_wdata),
       .m14_axi_wstrb(m14_axi_wstrb),
       .m14_axi_wlast(m14_axi_wlast),
       .m14_axi_bvalid(m14_axi_bvalid),
       .m14_axi_bready(m14_axi_bready),
       .m14_axi_arvalid(m14_axi_arvalid),
       .m14_axi_arready(m14_axi_arready),
       .m14_axi_araddr(m14_axi_araddr),
       .m14_axi_arlen(m14_axi_arlen),
       .m14_axi_rvalid(m14_axi_rvalid),
       .m14_axi_rready(m14_axi_rready),
       .m14_axi_rdata(m14_axi_rdata),
       .m14_axi_rlast(m14_axi_rlast),

       .m15_axi_awvalid(m15_axi_awvalid),
       .m15_axi_awready(m15_axi_awready),
       .m15_axi_awaddr(m15_axi_awaddr),
       .m15_axi_awlen(m15_axi_awlen),
       .m15_axi_wvalid(m15_axi_wvalid),
       .m15_axi_wready(m15_axi_wready),
       .m15_axi_wdata(m15_axi_wdata),
       .m15_axi_wstrb(m15_axi_wstrb),
       .m15_axi_wlast(m15_axi_wlast),
       .m15_axi_bvalid(m15_axi_bvalid),
       .m15_axi_bready(m15_axi_bready),
       .m15_axi_arvalid(m15_axi_arvalid),
       .m15_axi_arready(m15_axi_arready),
       .m15_axi_araddr(m15_axi_araddr),
       .m15_axi_arlen(m15_axi_arlen),
       .m15_axi_rvalid(m15_axi_rvalid),
       .m15_axi_rready(m15_axi_rready),
       .m15_axi_rdata(m15_axi_rdata),
       .m15_axi_rlast(m15_axi_rlast),

       .m16_axi_awvalid(m16_axi_awvalid),
       .m16_axi_awready(m16_axi_awready),
       .m16_axi_awaddr(m16_axi_awaddr),
       .m16_axi_awlen(m16_axi_awlen),
       .m16_axi_wvalid(m16_axi_wvalid),
       .m16_axi_wready(m16_axi_wready),
       .m16_axi_wdata(m16_axi_wdata),
       .m16_axi_wstrb(m16_axi_wstrb),
       .m16_axi_wlast(m16_axi_wlast),
       .m16_axi_bvalid(m16_axi_bvalid),
       .m16_axi_bready(m16_axi_bready),
       .m16_axi_arvalid(m16_axi_arvalid),
       .m16_axi_arready(m16_axi_arready),
       .m16_axi_araddr(m16_axi_araddr),
       .m16_axi_arlen(m16_axi_arlen),
       .m16_axi_rvalid(m16_axi_rvalid),
       .m16_axi_rready(m16_axi_rready),
       .m16_axi_rdata(m16_axi_rdata),
       .m16_axi_rlast(m16_axi_rlast),

       .m17_axi_awvalid(m17_axi_awvalid),
       .m17_axi_awready(m17_axi_awready),
       .m17_axi_awaddr(m17_axi_awaddr),
       .m17_axi_awlen(m17_axi_awlen),
       .m17_axi_wvalid(m17_axi_wvalid),
       .m17_axi_wready(m17_axi_wready),
       .m17_axi_wdata(m17_axi_wdata),
       .m17_axi_wstrb(m17_axi_wstrb),
       .m17_axi_wlast(m17_axi_wlast),
       .m17_axi_bvalid(m17_axi_bvalid),
       .m17_axi_bready(m17_axi_bready),
       .m17_axi_arvalid(m17_axi_arvalid),
       .m17_axi_arready(m17_axi_arready),
       .m17_axi_araddr(m17_axi_araddr),
       .m17_axi_arlen(m17_axi_arlen),
       .m17_axi_rvalid(m17_axi_rvalid),
       .m17_axi_rready(m17_axi_rready),
       .m17_axi_rdata(m17_axi_rdata),
       .m17_axi_rlast(m17_axi_rlast),

       .m18_axi_awvalid(m18_axi_awvalid),
       .m18_axi_awready(m18_axi_awready),
       .m18_axi_awaddr(m18_axi_awaddr),
       .m18_axi_awlen(m18_axi_awlen),
       .m18_axi_wvalid(m18_axi_wvalid),
       .m18_axi_wready(m18_axi_wready),
       .m18_axi_wdata(m18_axi_wdata),
       .m18_axi_wstrb(m18_axi_wstrb),
       .m18_axi_wlast(m18_axi_wlast),
       .m18_axi_bvalid(m18_axi_bvalid),
       .m18_axi_bready(m18_axi_bready),
       .m18_axi_arvalid(m18_axi_arvalid),
       .m18_axi_arready(m18_axi_arready),
       .m18_axi_araddr(m18_axi_araddr),
       .m18_axi_arlen(m18_axi_arlen),
       .m18_axi_rvalid(m18_axi_rvalid),
       .m18_axi_rready(m18_axi_rready),
       .m18_axi_rdata(m18_axi_rdata),
       .m18_axi_rlast(m18_axi_rlast),

       .m19_axi_awvalid(m19_axi_awvalid),
       .m19_axi_awready(m19_axi_awready),
       .m19_axi_awaddr(m19_axi_awaddr),
       .m19_axi_awlen(m19_axi_awlen),
       .m19_axi_wvalid(m19_axi_wvalid),
       .m19_axi_wready(m19_axi_wready),
       .m19_axi_wdata(m19_axi_wdata),
       .m19_axi_wstrb(m19_axi_wstrb),
       .m19_axi_wlast(m19_axi_wlast),
       .m19_axi_bvalid(m19_axi_bvalid),
       .m19_axi_bready(m19_axi_bready),
       .m19_axi_arvalid(m19_axi_arvalid),
       .m19_axi_arready(m19_axi_arready),
       .m19_axi_araddr(m19_axi_araddr),
       .m19_axi_arlen(m19_axi_arlen),
       .m19_axi_rvalid(m19_axi_rvalid),
       .m19_axi_rready(m19_axi_rready),
       .m19_axi_rdata(m19_axi_rdata),
       .m19_axi_rlast(m19_axi_rlast),

       .m20_axi_awvalid(m20_axi_awvalid),
       .m20_axi_awready(m20_axi_awready),
       .m20_axi_awaddr(m20_axi_awaddr),
       .m20_axi_awlen(m20_axi_awlen),
       .m20_axi_wvalid(m20_axi_wvalid),
       .m20_axi_wready(m20_axi_wready),
       .m20_axi_wdata(m20_axi_wdata),
       .m20_axi_wstrb(m20_axi_wstrb),
       .m20_axi_wlast(m20_axi_wlast),
       .m20_axi_bvalid(m20_axi_bvalid),
       .m20_axi_bready(m20_axi_bready),
       .m20_axi_arvalid(m20_axi_arvalid),
       .m20_axi_arready(m20_axi_arready),
       .m20_axi_araddr(m20_axi_araddr),
       .m20_axi_arlen(m20_axi_arlen),
       .m20_axi_rvalid(m20_axi_rvalid),
       .m20_axi_rready(m20_axi_rready),
       .m20_axi_rdata(m20_axi_rdata),
       .m20_axi_rlast(m20_axi_rlast),

       .m21_axi_awvalid(m21_axi_awvalid),
       .m21_axi_awready(m21_axi_awready),
       .m21_axi_awaddr(m21_axi_awaddr),
       .m21_axi_awlen(m21_axi_awlen),
       .m21_axi_wvalid(m21_axi_wvalid),
       .m21_axi_wready(m21_axi_wready),
       .m21_axi_wdata(m21_axi_wdata),
       .m21_axi_wstrb(m21_axi_wstrb),
       .m21_axi_wlast(m21_axi_wlast),
       .m21_axi_bvalid(m21_axi_bvalid),
       .m21_axi_bready(m21_axi_bready),
       .m21_axi_arvalid(m21_axi_arvalid),
       .m21_axi_arready(m21_axi_arready),
       .m21_axi_araddr(m21_axi_araddr),
       .m21_axi_arlen(m21_axi_arlen),
       .m21_axi_rvalid(m21_axi_rvalid),
       .m21_axi_rready(m21_axi_rready),
       .m21_axi_rdata(m21_axi_rdata),
       .m21_axi_rlast(m21_axi_rlast),

       .m22_axi_awvalid(m22_axi_awvalid),
       .m22_axi_awready(m22_axi_awready),
       .m22_axi_awaddr(m22_axi_awaddr),
       .m22_axi_awlen(m22_axi_awlen),
       .m22_axi_wvalid(m22_axi_wvalid),
       .m22_axi_wready(m22_axi_wready),
       .m22_axi_wdata(m22_axi_wdata),
       .m22_axi_wstrb(m22_axi_wstrb),
       .m22_axi_wlast(m22_axi_wlast),
       .m22_axi_bvalid(m22_axi_bvalid),
       .m22_axi_bready(m22_axi_bready),
       .m22_axi_arvalid(m22_axi_arvalid),
       .m22_axi_arready(m22_axi_arready),
       .m22_axi_araddr(m22_axi_araddr),
       .m22_axi_arlen(m22_axi_arlen),
       .m22_axi_rvalid(m22_axi_rvalid),
       .m22_axi_rready(m22_axi_rready),
       .m22_axi_rdata(m22_axi_rdata),
       .m22_axi_rlast(m22_axi_rlast),

       .m23_axi_awvalid(m23_axi_awvalid),
       .m23_axi_awready(m23_axi_awready),
       .m23_axi_awaddr(m23_axi_awaddr),
       .m23_axi_awlen(m23_axi_awlen),
       .m23_axi_wvalid(m23_axi_wvalid),
       .m23_axi_wready(m23_axi_wready),
       .m23_axi_wdata(m23_axi_wdata),
       .m23_axi_wstrb(m23_axi_wstrb),
       .m23_axi_wlast(m23_axi_wlast),
       .m23_axi_bvalid(m23_axi_bvalid),
       .m23_axi_bready(m23_axi_bready),
       .m23_axi_arvalid(m23_axi_arvalid),
       .m23_axi_arready(m23_axi_arready),
       .m23_axi_araddr(m23_axi_araddr),
       .m23_axi_arlen(m23_axi_arlen),
       .m23_axi_rvalid(m23_axi_rvalid),
       .m23_axi_rready(m23_axi_rready),
       .m23_axi_rdata(m23_axi_rdata),
       .m23_axi_rlast(m23_axi_rlast),

       .m24_axi_awvalid(m24_axi_awvalid),
       .m24_axi_awready(m24_axi_awready),
       .m24_axi_awaddr(m24_axi_awaddr),
       .m24_axi_awlen(m24_axi_awlen),
       .m24_axi_wvalid(m24_axi_wvalid),
       .m24_axi_wready(m24_axi_wready),
       .m24_axi_wdata(m24_axi_wdata),
       .m24_axi_wstrb(m24_axi_wstrb),
       .m24_axi_wlast(m24_axi_wlast),
       .m24_axi_bvalid(m24_axi_bvalid),
       .m24_axi_bready(m24_axi_bready),
       .m24_axi_arvalid(m24_axi_arvalid),
       .m24_axi_arready(m24_axi_arready),
       .m24_axi_araddr(m24_axi_araddr),
       .m24_axi_arlen(m24_axi_arlen),
       .m24_axi_rvalid(m24_axi_rvalid),
       .m24_axi_rready(m24_axi_rready),
       .m24_axi_rdata(m24_axi_rdata),
       .m24_axi_rlast(m24_axi_rlast),

       .m25_axi_awvalid(m25_axi_awvalid),
       .m25_axi_awready(m25_axi_awready),
       .m25_axi_awaddr(m25_axi_awaddr),
       .m25_axi_awlen(m25_axi_awlen),
       .m25_axi_wvalid(m25_axi_wvalid),
       .m25_axi_wready(m25_axi_wready),
       .m25_axi_wdata(m25_axi_wdata),
       .m25_axi_wstrb(m25_axi_wstrb),
       .m25_axi_wlast(m25_axi_wlast),
       .m25_axi_bvalid(m25_axi_bvalid),
       .m25_axi_bready(m25_axi_bready),
       .m25_axi_arvalid(m25_axi_arvalid),
       .m25_axi_arready(m25_axi_arready),
       .m25_axi_araddr(m25_axi_araddr),
       .m25_axi_arlen(m25_axi_arlen),
       .m25_axi_rvalid(m25_axi_rvalid),
       .m25_axi_rready(m25_axi_rready),
       .m25_axi_rdata(m25_axi_rdata),
       .m25_axi_rlast(m25_axi_rlast),

       .m26_axi_awvalid(m26_axi_awvalid),
       .m26_axi_awready(m26_axi_awready),
       .m26_axi_awaddr(m26_axi_awaddr),
       .m26_axi_awlen(m26_axi_awlen),
       .m26_axi_wvalid(m26_axi_wvalid),
       .m26_axi_wready(m26_axi_wready),
       .m26_axi_wdata(m26_axi_wdata),
       .m26_axi_wstrb(m26_axi_wstrb),
       .m26_axi_wlast(m26_axi_wlast),
       .m26_axi_bvalid(m26_axi_bvalid),
       .m26_axi_bready(m26_axi_bready),
       .m26_axi_arvalid(m26_axi_arvalid),
       .m26_axi_arready(m26_axi_arready),
       .m26_axi_araddr(m26_axi_araddr),
       .m26_axi_arlen(m26_axi_arlen),
       .m26_axi_rvalid(m26_axi_rvalid),
       .m26_axi_rready(m26_axi_rready),
       .m26_axi_rdata(m26_axi_rdata),
       .m26_axi_rlast(m26_axi_rlast),

       .m27_axi_awvalid(m27_axi_awvalid),
       .m27_axi_awready(m27_axi_awready),
       .m27_axi_awaddr(m27_axi_awaddr),
       .m27_axi_awlen(m27_axi_awlen),
       .m27_axi_wvalid(m27_axi_wvalid),
       .m27_axi_wready(m27_axi_wready),
       .m27_axi_wdata(m27_axi_wdata),
       .m27_axi_wstrb(m27_axi_wstrb),
       .m27_axi_wlast(m27_axi_wlast),
       .m27_axi_bvalid(m27_axi_bvalid),
       .m27_axi_bready(m27_axi_bready),
       .m27_axi_arvalid(m27_axi_arvalid),
       .m27_axi_arready(m27_axi_arready),
       .m27_axi_araddr(m27_axi_araddr),
       .m27_axi_arlen(m27_axi_arlen),
       .m27_axi_rvalid(m27_axi_rvalid),
       .m27_axi_rready(m27_axi_rready),
       .m27_axi_rdata(m27_axi_rdata),
       .m27_axi_rlast(m27_axi_rlast),

       .m28_axi_awvalid(m28_axi_awvalid),
       .m28_axi_awready(m28_axi_awready),
       .m28_axi_awaddr(m28_axi_awaddr),
       .m28_axi_awlen(m28_axi_awlen),
       .m28_axi_wvalid(m28_axi_wvalid),
       .m28_axi_wready(m28_axi_wready),
       .m28_axi_wdata(m28_axi_wdata),
       .m28_axi_wstrb(m28_axi_wstrb),
       .m28_axi_wlast(m28_axi_wlast),
       .m28_axi_bvalid(m28_axi_bvalid),
       .m28_axi_bready(m28_axi_bready),
       .m28_axi_arvalid(m28_axi_arvalid),
       .m28_axi_arready(m28_axi_arready),
       .m28_axi_araddr(m28_axi_araddr),
       .m28_axi_arlen(m28_axi_arlen),
       .m28_axi_rvalid(m28_axi_rvalid),
       .m28_axi_rready(m28_axi_rready),
       .m28_axi_rdata(m28_axi_rdata),
       .m28_axi_rlast(m28_axi_rlast),

       .m29_axi_awvalid(m29_axi_awvalid),
       .m29_axi_awready(m29_axi_awready),
       .m29_axi_awaddr(m29_axi_awaddr),
       .m29_axi_awlen(m29_axi_awlen),
       .m29_axi_wvalid(m29_axi_wvalid),
       .m29_axi_wready(m29_axi_wready),
       .m29_axi_wdata(m29_axi_wdata),
       .m29_axi_wstrb(m29_axi_wstrb),
       .m29_axi_wlast(m29_axi_wlast),
       .m29_axi_bvalid(m29_axi_bvalid),
       .m29_axi_bready(m29_axi_bready),
       .m29_axi_arvalid(m29_axi_arvalid),
       .m29_axi_arready(m29_axi_arready),
       .m29_axi_araddr(m29_axi_araddr),
       .m29_axi_arlen(m29_axi_arlen),
       .m29_axi_rvalid(m29_axi_rvalid),
       .m29_axi_rready(m29_axi_rready),
       .m29_axi_rdata(m29_axi_rdata),
       .m29_axi_rlast(m29_axi_rlast),

       .m30_axi_awvalid(m30_axi_awvalid),
       .m30_axi_awready(m30_axi_awready),
       .m30_axi_awaddr(m30_axi_awaddr),
       .m30_axi_awlen(m30_axi_awlen),
       .m30_axi_wvalid(m30_axi_wvalid),
       .m30_axi_wready(m30_axi_wready),
       .m30_axi_wdata(m30_axi_wdata),
       .m30_axi_wstrb(m30_axi_wstrb),
       .m30_axi_wlast(m30_axi_wlast),
       .m30_axi_bvalid(m30_axi_bvalid),
       .m30_axi_bready(m30_axi_bready),
       .m30_axi_arvalid(m30_axi_arvalid),
       .m30_axi_arready(m30_axi_arready),
       .m30_axi_araddr(m30_axi_araddr),
       .m30_axi_arlen(m30_axi_arlen),
       .m30_axi_rvalid(m30_axi_rvalid),
       .m30_axi_rready(m30_axi_rready),
       .m30_axi_rdata(m30_axi_rdata),
       .m30_axi_rlast(m30_axi_rlast),

       .m31_axi_awvalid(m31_axi_awvalid),
       .m31_axi_awready(m31_axi_awready),
       .m31_axi_awaddr(m31_axi_awaddr),
       .m31_axi_awlen(m31_axi_awlen),
       .m31_axi_wvalid(m31_axi_wvalid),
       .m31_axi_wready(m31_axi_wready),
       .m31_axi_wdata(m31_axi_wdata),
       .m31_axi_wstrb(m31_axi_wstrb),
       .m31_axi_wlast(m31_axi_wlast),
       .m31_axi_bvalid(m31_axi_bvalid),
       .m31_axi_bready(m31_axi_bready),
       .m31_axi_arvalid(m31_axi_arvalid),
       .m31_axi_arready(m31_axi_arready),
       .m31_axi_araddr(m31_axi_araddr),
       .m31_axi_arlen(m31_axi_arlen),
       .m31_axi_rvalid(m31_axi_rvalid),
       .m31_axi_rready(m31_axi_rready),
       .m31_axi_rdata(m31_axi_rdata),
       .m31_axi_rlast(m31_axi_rlast),

       .s_axi_control_awvalid(s_axi_control_awvalid),
       .s_axi_control_awready(s_axi_control_awready),
       .s_axi_control_awaddr(s_axi_control_awaddr),
       .s_axi_control_wvalid(s_axi_control_wvalid),
       .s_axi_control_wready(s_axi_control_wready),
       .s_axi_control_wdata(s_axi_control_wdata),
       .s_axi_control_wstrb(s_axi_control_wstrb),
       .s_axi_control_arvalid(s_axi_control_arvalid),
       .s_axi_control_arready(s_axi_control_arready),
       .s_axi_control_araddr(s_axi_control_araddr),
       .s_axi_control_rvalid(s_axi_control_rvalid),
       .s_axi_control_rready(s_axi_control_rready),
       .s_axi_control_rdata(s_axi_control_rdata),
       .s_axi_control_rresp(s_axi_control_rresp),
       .s_axi_control_bvalid(s_axi_control_bvalid),
       .s_axi_control_bready(s_axi_control_bready),
       .s_axi_control_bresp(s_axi_control_bresp),

       .interrupt(interrupt)
       );

endmodule
